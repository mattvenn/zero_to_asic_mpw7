magic
tech sky130B
magscale 1 2
timestamp 1661721994
<< obsli1 >>
rect 0 0 584000 704000
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 37182 702788 37188 702840
rect 37240 702828 37246 702840
rect 202782 702828 202788 702840
rect 37240 702800 202788 702828
rect 37240 702788 37246 702800
rect 202782 702788 202788 702800
rect 202840 702788 202846 702840
rect 63402 702720 63408 702772
rect 63460 702760 63466 702772
rect 267642 702760 267648 702772
rect 63460 702732 267648 702760
rect 63460 702720 63466 702732
rect 267642 702720 267648 702732
rect 267700 702720 267706 702772
rect 297358 702720 297364 702772
rect 297416 702760 297422 702772
rect 494790 702760 494796 702772
rect 297416 702732 494796 702760
rect 297416 702720 297422 702732
rect 494790 702720 494796 702732
rect 494848 702720 494854 702772
rect 8110 702652 8116 702704
rect 8168 702692 8174 702704
rect 210418 702692 210424 702704
rect 8168 702664 210424 702692
rect 8168 702652 8174 702664
rect 210418 702652 210424 702664
rect 210476 702652 210482 702704
rect 248322 702652 248328 702704
rect 248380 702692 248386 702704
rect 527174 702692 527180 702704
rect 248380 702664 527180 702692
rect 248380 702652 248386 702664
rect 527174 702652 527180 702664
rect 527232 702652 527238 702704
rect 130378 702584 130384 702636
rect 130436 702624 130442 702636
rect 413646 702624 413652 702636
rect 130436 702596 413652 702624
rect 130436 702584 130442 702596
rect 413646 702584 413652 702596
rect 413704 702584 413710 702636
rect 53742 702516 53748 702568
rect 53800 702556 53806 702568
rect 462314 702556 462320 702568
rect 53800 702528 462320 702556
rect 53800 702516 53806 702528
rect 462314 702516 462320 702528
rect 462372 702516 462378 702568
rect 63310 702448 63316 702500
rect 63368 702488 63374 702500
rect 543458 702488 543464 702500
rect 63368 702460 543464 702488
rect 63368 702448 63374 702460
rect 543458 702448 543464 702460
rect 543516 702448 543522 702500
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 48958 700380 48964 700392
rect 24360 700352 48964 700380
rect 24360 700340 24366 700352
rect 48958 700340 48964 700352
rect 49016 700340 49022 700392
rect 45462 700272 45468 700324
rect 45520 700312 45526 700324
rect 137830 700312 137836 700324
rect 45520 700284 137836 700312
rect 45520 700272 45526 700284
rect 137830 700272 137836 700284
rect 137888 700272 137894 700324
rect 235166 700272 235172 700324
rect 235224 700312 235230 700324
rect 244274 700312 244280 700324
rect 235224 700284 244280 700312
rect 235224 700272 235230 700284
rect 244274 700272 244280 700284
rect 244332 700272 244338 700324
rect 253198 700272 253204 700324
rect 253256 700312 253262 700324
rect 559650 700312 559656 700324
rect 253256 700284 559656 700312
rect 253256 700272 253262 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 100018 699660 100024 699712
rect 100076 699700 100082 699712
rect 105446 699700 105452 699712
rect 100076 699672 105452 699700
rect 100076 699660 100082 699672
rect 105446 699660 105452 699672
rect 105504 699660 105510 699712
rect 395338 699660 395344 699712
rect 395396 699700 395402 699712
rect 397454 699700 397460 699712
rect 395396 699672 397460 699700
rect 395396 699660 395402 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 63494 698912 63500 698964
rect 63552 698952 63558 698964
rect 218974 698952 218980 698964
rect 63552 698924 218980 698952
rect 63552 698912 63558 698924
rect 218974 698912 218980 698924
rect 219032 698912 219038 698964
rect 262122 698912 262128 698964
rect 262180 698952 262186 698964
rect 429838 698952 429844 698964
rect 262180 698924 429844 698952
rect 262180 698912 262186 698924
rect 429838 698912 429844 698924
rect 429896 698912 429902 698964
rect 278038 697552 278044 697604
rect 278096 697592 278102 697604
rect 348786 697592 348792 697604
rect 278096 697564 348792 697592
rect 278096 697552 278102 697564
rect 348786 697552 348792 697564
rect 348844 697552 348850 697604
rect 363598 696940 363604 696992
rect 363656 696980 363662 696992
rect 580166 696980 580172 696992
rect 363656 696952 580172 696980
rect 363656 696940 363662 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 46198 683176 46204 683188
rect 3476 683148 46204 683176
rect 3476 683136 3482 683148
rect 46198 683136 46204 683148
rect 46256 683136 46262 683188
rect 242802 683136 242808 683188
rect 242860 683176 242866 683188
rect 580166 683176 580172 683188
rect 242860 683148 580172 683176
rect 242860 683136 242866 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 291838 670692 291844 670744
rect 291896 670732 291902 670744
rect 580166 670732 580172 670744
rect 291896 670704 580172 670732
rect 291896 670692 291902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 43438 656928 43444 656940
rect 3568 656900 43444 656928
rect 3568 656888 3574 656900
rect 43438 656888 43444 656900
rect 43496 656888 43502 656940
rect 251082 643084 251088 643136
rect 251140 643124 251146 643136
rect 580166 643124 580172 643136
rect 251140 643096 580172 643124
rect 251140 643084 251146 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 229738 632108 229744 632120
rect 3568 632080 229744 632108
rect 3568 632068 3574 632080
rect 229738 632068 229744 632080
rect 229796 632068 229802 632120
rect 175366 630640 175372 630692
rect 175424 630680 175430 630692
rect 244366 630680 244372 630692
rect 175424 630652 244372 630680
rect 175424 630640 175430 630652
rect 244366 630640 244372 630652
rect 244424 630680 244430 630692
rect 580166 630680 580172 630692
rect 244424 630652 580172 630680
rect 244424 630640 244430 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 618604 3516 618656
rect 3568 618644 3574 618656
rect 7558 618644 7564 618656
rect 3568 618616 7564 618644
rect 3568 618604 3574 618616
rect 7558 618604 7564 618616
rect 7616 618604 7622 618656
rect 48958 607112 48964 607164
rect 49016 607152 49022 607164
rect 52270 607152 52276 607164
rect 49016 607124 52276 607152
rect 49016 607112 49022 607124
rect 52270 607112 52276 607124
rect 52328 607112 52334 607164
rect 3510 606024 3516 606076
rect 3568 606064 3574 606076
rect 8938 606064 8944 606076
rect 3568 606036 8944 606064
rect 3568 606024 3574 606036
rect 8938 606024 8944 606036
rect 8996 606024 9002 606076
rect 52270 605820 52276 605872
rect 52328 605860 52334 605872
rect 185026 605860 185032 605872
rect 52328 605832 185032 605860
rect 52328 605820 52334 605832
rect 185026 605820 185032 605832
rect 185084 605820 185090 605872
rect 88334 600924 88340 600976
rect 88392 600964 88398 600976
rect 236638 600964 236644 600976
rect 88392 600936 236644 600964
rect 88392 600924 88398 600936
rect 236638 600924 236644 600936
rect 236696 600924 236702 600976
rect 71774 599564 71780 599616
rect 71832 599604 71838 599616
rect 245746 599604 245752 599616
rect 71832 599576 245752 599604
rect 71832 599564 71838 599576
rect 245746 599564 245752 599576
rect 245804 599564 245810 599616
rect 40034 596776 40040 596828
rect 40092 596816 40098 596828
rect 217318 596816 217324 596828
rect 40092 596788 217324 596816
rect 40092 596776 40098 596788
rect 217318 596776 217324 596788
rect 217376 596776 217382 596828
rect 169754 595416 169760 595468
rect 169812 595456 169818 595468
rect 245838 595456 245844 595468
rect 169812 595428 245844 595456
rect 169812 595416 169818 595428
rect 245838 595416 245844 595428
rect 245896 595416 245902 595468
rect 3418 594056 3424 594108
rect 3476 594096 3482 594108
rect 244550 594096 244556 594108
rect 3476 594068 244556 594096
rect 3476 594056 3482 594068
rect 244550 594056 244556 594068
rect 244608 594056 244614 594108
rect 256602 594056 256608 594108
rect 256660 594096 256666 594108
rect 299474 594096 299480 594108
rect 256660 594068 299480 594096
rect 256660 594056 256666 594068
rect 299474 594056 299480 594068
rect 299532 594056 299538 594108
rect 90174 592628 90180 592680
rect 90232 592668 90238 592680
rect 100018 592668 100024 592680
rect 90232 592640 100024 592668
rect 90232 592628 90238 592640
rect 100018 592628 100024 592640
rect 100076 592628 100082 592680
rect 220722 592628 220728 592680
rect 220780 592668 220786 592680
rect 282914 592668 282920 592680
rect 220780 592640 282920 592668
rect 220780 592628 220786 592640
rect 282914 592628 282920 592640
rect 282972 592628 282978 592680
rect 46842 592152 46848 592204
rect 46900 592192 46906 592204
rect 102594 592192 102600 592204
rect 46900 592164 102600 592192
rect 46900 592152 46906 592164
rect 102594 592152 102600 592164
rect 102652 592152 102658 592204
rect 45278 592084 45284 592136
rect 45336 592124 45342 592136
rect 134150 592124 134156 592136
rect 45336 592096 134156 592124
rect 45336 592084 45342 592096
rect 134150 592084 134156 592096
rect 134208 592084 134214 592136
rect 48130 592016 48136 592068
rect 48188 592056 48194 592068
rect 153470 592056 153476 592068
rect 48188 592028 153476 592056
rect 48188 592016 48194 592028
rect 153470 592016 153476 592028
rect 153528 592016 153534 592068
rect 153194 591268 153200 591320
rect 153252 591308 153258 591320
rect 251174 591308 251180 591320
rect 153252 591280 251180 591308
rect 153252 591268 153258 591280
rect 251174 591268 251180 591280
rect 251232 591268 251238 591320
rect 53650 590860 53656 590912
rect 53708 590900 53714 590912
rect 86494 590900 86500 590912
rect 53708 590872 86500 590900
rect 53708 590860 53714 590872
rect 86494 590860 86500 590872
rect 86552 590860 86558 590912
rect 42610 590792 42616 590844
rect 42668 590832 42674 590844
rect 112254 590832 112260 590844
rect 42668 590804 112260 590832
rect 42668 590792 42674 590804
rect 112254 590792 112260 590804
rect 112312 590792 112318 590844
rect 44082 590724 44088 590776
rect 44140 590764 44146 590776
rect 143810 590764 143816 590776
rect 44140 590736 143816 590764
rect 44140 590724 44146 590736
rect 143810 590724 143816 590736
rect 143868 590724 143874 590776
rect 46750 590656 46756 590708
rect 46808 590696 46814 590708
rect 159910 590696 159916 590708
rect 46808 590668 159916 590696
rect 46808 590656 46814 590668
rect 159910 590656 159916 590668
rect 159968 590656 159974 590708
rect 130378 590248 130384 590300
rect 130436 590288 130442 590300
rect 130930 590288 130936 590300
rect 130436 590260 130936 590288
rect 130436 590248 130442 590260
rect 130930 590248 130936 590260
rect 130988 590248 130994 590300
rect 201402 589908 201408 589960
rect 201460 589948 201466 589960
rect 580166 589948 580172 589960
rect 201460 589920 580172 589948
rect 201460 589908 201466 589920
rect 580166 589908 580172 589920
rect 580224 589908 580230 589960
rect 55030 589636 55036 589688
rect 55088 589676 55094 589688
rect 118694 589676 118700 589688
rect 55088 589648 118700 589676
rect 55088 589636 55094 589648
rect 118694 589636 118700 589648
rect 118752 589636 118758 589688
rect 53558 589568 53564 589620
rect 53616 589608 53622 589620
rect 121914 589608 121920 589620
rect 53616 589580 121920 589608
rect 53616 589568 53622 589580
rect 121914 589568 121920 589580
rect 121972 589568 121978 589620
rect 61930 589500 61936 589552
rect 61988 589540 61994 589552
rect 130930 589540 130936 589552
rect 61988 589512 130936 589540
rect 61988 589500 61994 589512
rect 130930 589500 130936 589512
rect 130988 589500 130994 589552
rect 52178 589432 52184 589484
rect 52236 589472 52242 589484
rect 140590 589472 140596 589484
rect 52236 589444 140596 589472
rect 52236 589432 52242 589444
rect 140590 589432 140596 589444
rect 140648 589432 140654 589484
rect 42702 589364 42708 589416
rect 42760 589404 42766 589416
rect 156690 589404 156696 589416
rect 42760 589376 156696 589404
rect 42760 589364 42766 589376
rect 156690 589364 156696 589376
rect 156748 589364 156754 589416
rect 35802 589296 35808 589348
rect 35860 589336 35866 589348
rect 163130 589336 163136 589348
rect 35860 589308 163136 589336
rect 35860 589296 35866 589308
rect 163130 589296 163136 589308
rect 163188 589296 163194 589348
rect 235994 589296 236000 589348
rect 236052 589336 236058 589348
rect 236638 589336 236644 589348
rect 236052 589308 236644 589336
rect 236052 589296 236058 589308
rect 236638 589296 236644 589308
rect 236696 589336 236702 589348
rect 258074 589336 258080 589348
rect 236696 589308 258080 589336
rect 236696 589296 236702 589308
rect 258074 589296 258080 589308
rect 258132 589296 258138 589348
rect 256694 588548 256700 588600
rect 256752 588588 256758 588600
rect 331214 588588 331220 588600
rect 256752 588560 331220 588588
rect 256752 588548 256758 588560
rect 331214 588548 331220 588560
rect 331272 588548 331278 588600
rect 56410 588208 56416 588260
rect 56468 588248 56474 588260
rect 90174 588248 90180 588260
rect 56468 588220 90180 588248
rect 56468 588208 56474 588220
rect 90174 588208 90180 588220
rect 90232 588208 90238 588260
rect 39666 588140 39672 588192
rect 39724 588180 39730 588192
rect 105906 588180 105912 588192
rect 39724 588152 105912 588180
rect 39724 588140 39730 588152
rect 105906 588140 105912 588152
rect 105964 588140 105970 588192
rect 229738 588140 229744 588192
rect 229796 588180 229802 588192
rect 249794 588180 249800 588192
rect 229796 588152 249800 588180
rect 229796 588140 229802 588152
rect 249794 588140 249800 588152
rect 249852 588140 249858 588192
rect 60090 588072 60096 588124
rect 60148 588112 60154 588124
rect 127802 588112 127808 588124
rect 60148 588084 127808 588112
rect 60148 588072 60154 588084
rect 127802 588072 127808 588084
rect 127860 588072 127866 588124
rect 226334 588072 226340 588124
rect 226392 588112 226398 588124
rect 256694 588112 256700 588124
rect 226392 588084 256700 588112
rect 226392 588072 226398 588084
rect 256694 588072 256700 588084
rect 256752 588072 256758 588124
rect 54938 588004 54944 588056
rect 54996 588044 55002 588056
rect 191558 588044 191564 588056
rect 54996 588016 191564 588044
rect 54996 588004 55002 588016
rect 191558 588004 191564 588016
rect 191616 588004 191622 588056
rect 210418 588004 210424 588056
rect 210476 588044 210482 588056
rect 244458 588044 244464 588056
rect 210476 588016 244464 588044
rect 210476 588004 210482 588016
rect 244458 588004 244464 588016
rect 244516 588004 244522 588056
rect 5442 587936 5448 587988
rect 5500 587976 5506 587988
rect 147122 587976 147128 587988
rect 5500 587948 147128 587976
rect 5500 587936 5506 587948
rect 147122 587936 147128 587948
rect 147180 587936 147186 587988
rect 242802 587936 242808 587988
rect 242860 587976 242866 587988
rect 289078 587976 289084 587988
rect 242860 587948 289084 587976
rect 242860 587936 242866 587948
rect 289078 587936 289084 587948
rect 289136 587936 289142 587988
rect 48958 587868 48964 587920
rect 49016 587908 49022 587920
rect 197998 587908 198004 587920
rect 49016 587880 198004 587908
rect 49016 587868 49022 587880
rect 197998 587868 198004 587880
rect 198056 587908 198062 587920
rect 246298 587908 246304 587920
rect 198056 587880 246304 587908
rect 198056 587868 198062 587880
rect 246298 587868 246304 587880
rect 246356 587868 246362 587920
rect 35158 586916 35164 586968
rect 35216 586956 35222 586968
rect 80146 586956 80152 586968
rect 35216 586928 80152 586956
rect 35216 586916 35222 586928
rect 80146 586916 80152 586928
rect 80204 586916 80210 586968
rect 34422 586848 34428 586900
rect 34480 586888 34486 586900
rect 77570 586888 77576 586900
rect 34480 586860 77576 586888
rect 34480 586848 34486 586860
rect 77570 586848 77576 586860
rect 77628 586848 77634 586900
rect 239214 586848 239220 586900
rect 239272 586888 239278 586900
rect 252554 586888 252560 586900
rect 239272 586860 252560 586888
rect 239272 586848 239278 586860
rect 252554 586848 252560 586860
rect 252612 586848 252618 586900
rect 49510 586780 49516 586832
rect 49568 586820 49574 586832
rect 96246 586820 96252 586832
rect 49568 586792 96252 586820
rect 49568 586780 49574 586792
rect 96246 586780 96252 586792
rect 96304 586780 96310 586832
rect 217318 586780 217324 586832
rect 217376 586820 217382 586832
rect 243170 586820 243176 586832
rect 217376 586792 243176 586820
rect 217376 586780 217382 586792
rect 243170 586780 243176 586792
rect 243228 586780 243234 586832
rect 59998 586712 60004 586764
rect 60056 586752 60062 586764
rect 109126 586752 109132 586764
rect 60056 586724 109132 586752
rect 60056 586712 60062 586724
rect 109126 586712 109132 586724
rect 109184 586712 109190 586764
rect 214098 586712 214104 586764
rect 214156 586752 214162 586764
rect 248414 586752 248420 586764
rect 214156 586724 248420 586752
rect 214156 586712 214162 586724
rect 248414 586712 248420 586724
rect 248472 586712 248478 586764
rect 62758 586644 62764 586696
rect 62816 586684 62822 586696
rect 115566 586684 115572 586696
rect 62816 586656 115572 586684
rect 62816 586644 62822 586656
rect 115566 586644 115572 586656
rect 115624 586644 115630 586696
rect 207658 586644 207664 586696
rect 207716 586684 207722 586696
rect 255314 586684 255320 586696
rect 207716 586656 255320 586684
rect 207716 586644 207722 586656
rect 255314 586644 255320 586656
rect 255372 586644 255378 586696
rect 79410 586576 79416 586628
rect 79468 586616 79474 586628
rect 137462 586616 137468 586628
rect 79468 586588 137468 586616
rect 79468 586576 79474 586588
rect 137462 586576 137468 586588
rect 137520 586576 137526 586628
rect 181898 586576 181904 586628
rect 181956 586616 181962 586628
rect 242986 586616 242992 586628
rect 181956 586588 242992 586616
rect 181956 586576 181962 586588
rect 242986 586576 242992 586588
rect 243044 586576 243050 586628
rect 63586 586508 63592 586560
rect 63644 586548 63650 586560
rect 150342 586548 150348 586560
rect 63644 586520 150348 586548
rect 63644 586508 63650 586520
rect 150342 586508 150348 586520
rect 150400 586508 150406 586560
rect 172882 586508 172888 586560
rect 172940 586548 172946 586560
rect 259454 586548 259460 586560
rect 172940 586520 259460 586548
rect 172940 586508 172946 586520
rect 259454 586508 259460 586520
rect 259512 586508 259518 586560
rect 63218 585760 63224 585812
rect 63276 585800 63282 585812
rect 79410 585800 79416 585812
rect 63276 585772 79416 585800
rect 63276 585760 63282 585772
rect 79410 585760 79416 585772
rect 79468 585760 79474 585812
rect 44818 585420 44824 585472
rect 44876 585460 44882 585472
rect 71130 585460 71136 585472
rect 44876 585432 71136 585460
rect 44876 585420 44882 585432
rect 71130 585420 71136 585432
rect 71188 585420 71194 585472
rect 41230 585352 41236 585404
rect 41288 585392 41294 585404
rect 67910 585392 67916 585404
rect 41288 585364 67916 585392
rect 41288 585352 41294 585364
rect 67910 585352 67916 585364
rect 67968 585352 67974 585404
rect 194778 585352 194784 585404
rect 194836 585392 194842 585404
rect 243630 585392 243636 585404
rect 194836 585364 243636 585392
rect 194836 585352 194842 585364
rect 243630 585352 243636 585364
rect 243688 585392 243694 585404
rect 251910 585392 251916 585404
rect 243688 585364 251916 585392
rect 243688 585352 243694 585364
rect 251910 585352 251916 585364
rect 251968 585352 251974 585404
rect 50338 585284 50344 585336
rect 50396 585324 50402 585336
rect 172882 585324 172888 585336
rect 50396 585296 172888 585324
rect 50396 585284 50402 585296
rect 172882 585284 172888 585296
rect 172940 585284 172946 585336
rect 220538 585284 220544 585336
rect 220596 585324 220602 585336
rect 220722 585324 220728 585336
rect 220596 585296 220728 585324
rect 220596 585284 220602 585296
rect 220722 585284 220728 585296
rect 220780 585324 220786 585336
rect 292574 585324 292580 585336
rect 220780 585296 292580 585324
rect 220780 585284 220786 585296
rect 292574 585284 292580 585296
rect 292632 585284 292638 585336
rect 31018 585216 31024 585268
rect 31076 585256 31082 585268
rect 263686 585256 263692 585268
rect 31076 585228 263692 585256
rect 31076 585216 31082 585228
rect 263686 585216 263692 585228
rect 263744 585216 263750 585268
rect 52362 585148 52368 585200
rect 52420 585188 52426 585200
rect 125226 585188 125232 585200
rect 52420 585160 125232 585188
rect 52420 585148 52426 585160
rect 125226 585148 125232 585160
rect 125284 585148 125290 585200
rect 166442 585148 166448 585200
rect 166500 585188 166506 585200
rect 245654 585188 245660 585200
rect 166500 585160 245660 585188
rect 166500 585148 166506 585160
rect 245654 585148 245660 585160
rect 245712 585148 245718 585200
rect 73982 584576 73988 584588
rect 64846 584548 73988 584576
rect 57882 583856 57888 583908
rect 57940 583896 57946 583908
rect 63586 583896 63592 583908
rect 57940 583868 63592 583896
rect 57940 583856 57946 583868
rect 63586 583856 63592 583868
rect 63644 583856 63650 583908
rect 49602 583788 49608 583840
rect 49660 583828 49666 583840
rect 64846 583828 64874 584548
rect 73982 584536 73988 584548
rect 74040 584536 74046 584588
rect 204714 584536 204720 584588
rect 204772 584576 204778 584588
rect 204772 584548 209774 584576
rect 204772 584536 204778 584548
rect 49660 583800 64874 583828
rect 209746 583828 209774 584548
rect 251266 583828 251272 583840
rect 209746 583800 251272 583828
rect 49660 583788 49666 583800
rect 251266 583788 251272 583800
rect 251324 583788 251330 583840
rect 2866 583720 2872 583772
rect 2924 583760 2930 583772
rect 57698 583760 57704 583772
rect 2924 583732 57704 583760
rect 2924 583720 2930 583732
rect 57698 583720 57704 583732
rect 57756 583760 57762 583772
rect 57882 583760 57888 583772
rect 57756 583732 57888 583760
rect 57756 583720 57762 583732
rect 57882 583720 57888 583732
rect 57940 583720 57946 583772
rect 58710 583720 58716 583772
rect 58768 583760 58774 583772
rect 247126 583760 247132 583772
rect 58768 583732 247132 583760
rect 58768 583720 58774 583732
rect 247126 583720 247132 583732
rect 247184 583720 247190 583772
rect 245654 582360 245660 582412
rect 245712 582400 245718 582412
rect 336734 582400 336740 582412
rect 245712 582372 336740 582400
rect 245712 582360 245718 582372
rect 336734 582360 336740 582372
rect 336792 582360 336798 582412
rect 243170 581612 243176 581664
rect 243228 581652 243234 581664
rect 276014 581652 276020 581664
rect 243228 581624 276020 581652
rect 243228 581612 243234 581624
rect 276014 581612 276020 581624
rect 276072 581612 276078 581664
rect 243262 578144 243268 578196
rect 243320 578184 243326 578196
rect 579798 578184 579804 578196
rect 243320 578156 579804 578184
rect 243320 578144 243326 578156
rect 579798 578144 579804 578156
rect 579856 578144 579862 578196
rect 245746 576512 245752 576564
rect 245804 576552 245810 576564
rect 245930 576552 245936 576564
rect 245804 576524 245936 576552
rect 245804 576512 245810 576524
rect 245930 576512 245936 576524
rect 245988 576512 245994 576564
rect 245746 575492 245752 575544
rect 245804 575532 245810 575544
rect 335354 575532 335360 575544
rect 245804 575504 335360 575532
rect 245804 575492 245810 575504
rect 335354 575492 335360 575504
rect 335412 575492 335418 575544
rect 245746 572704 245752 572756
rect 245804 572744 245810 572756
rect 287698 572744 287704 572756
rect 245804 572716 287704 572744
rect 245804 572704 245810 572716
rect 287698 572704 287704 572716
rect 287756 572704 287762 572756
rect 55122 568556 55128 568608
rect 55180 568596 55186 568608
rect 60734 568596 60740 568608
rect 55180 568568 60740 568596
rect 55180 568556 55186 568568
rect 60734 568556 60740 568568
rect 60792 568556 60798 568608
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 14458 565876 14464 565888
rect 3476 565848 14464 565876
rect 3476 565836 3482 565848
rect 14458 565836 14464 565848
rect 14516 565836 14522 565888
rect 245746 565836 245752 565888
rect 245804 565876 245810 565888
rect 332594 565876 332600 565888
rect 245804 565848 332600 565876
rect 245804 565836 245810 565848
rect 332594 565836 332600 565848
rect 332652 565836 332658 565888
rect 27522 564408 27528 564460
rect 27580 564448 27586 564460
rect 60734 564448 60740 564460
rect 27580 564420 60740 564448
rect 27580 564408 27586 564420
rect 60734 564408 60740 564420
rect 60792 564408 60798 564460
rect 445018 563048 445024 563100
rect 445076 563088 445082 563100
rect 580166 563088 580172 563100
rect 445076 563060 580172 563088
rect 445076 563048 445082 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 48222 561688 48228 561740
rect 48280 561728 48286 561740
rect 60734 561728 60740 561740
rect 48280 561700 60740 561728
rect 48280 561688 48286 561700
rect 60734 561688 60740 561700
rect 60792 561688 60798 561740
rect 245746 558900 245752 558952
rect 245804 558940 245810 558952
rect 248506 558940 248512 558952
rect 245804 558912 248512 558940
rect 245804 558900 245810 558912
rect 248506 558900 248512 558912
rect 248564 558900 248570 558952
rect 245746 556180 245752 556232
rect 245804 556220 245810 556232
rect 314654 556220 314660 556232
rect 245804 556192 314660 556220
rect 245804 556180 245810 556192
rect 314654 556180 314660 556192
rect 314712 556220 314718 556232
rect 500218 556220 500224 556232
rect 314712 556192 500224 556220
rect 314712 556180 314718 556192
rect 500218 556180 500224 556192
rect 500276 556180 500282 556232
rect 33042 554752 33048 554804
rect 33100 554792 33106 554804
rect 60734 554792 60740 554804
rect 33100 554764 60740 554792
rect 33100 554752 33106 554764
rect 60734 554752 60740 554764
rect 60792 554752 60798 554804
rect 3142 554684 3148 554736
rect 3200 554724 3206 554736
rect 31018 554724 31024 554736
rect 3200 554696 31024 554724
rect 3200 554684 3206 554696
rect 31018 554684 31024 554696
rect 31076 554684 31082 554736
rect 39850 552032 39856 552084
rect 39908 552072 39914 552084
rect 60734 552072 60740 552084
rect 39908 552044 60740 552072
rect 39908 552032 39914 552044
rect 60734 552032 60740 552044
rect 60792 552032 60798 552084
rect 264974 549856 264980 549908
rect 265032 549896 265038 549908
rect 363598 549896 363604 549908
rect 265032 549868 363604 549896
rect 265032 549856 265038 549868
rect 363598 549856 363604 549868
rect 363656 549856 363662 549908
rect 245746 549244 245752 549296
rect 245804 549284 245810 549296
rect 264974 549284 264980 549296
rect 245804 549256 264980 549284
rect 245804 549244 245810 549256
rect 264974 549244 264980 549256
rect 265032 549244 265038 549296
rect 57882 548360 57888 548412
rect 57940 548400 57946 548412
rect 60734 548400 60740 548412
rect 57940 548372 60740 548400
rect 57940 548360 57946 548372
rect 60734 548360 60740 548372
rect 60792 548360 60798 548412
rect 7558 542988 7564 543040
rect 7616 543028 7622 543040
rect 39942 543028 39948 543040
rect 7616 543000 39948 543028
rect 7616 542988 7622 543000
rect 39942 542988 39948 543000
rect 40000 542988 40006 543040
rect 39942 542376 39948 542428
rect 40000 542416 40006 542428
rect 60734 542416 60740 542428
rect 40000 542388 60740 542416
rect 40000 542376 40006 542388
rect 60734 542376 60740 542388
rect 60792 542376 60798 542428
rect 245746 539588 245752 539640
rect 245804 539628 245810 539640
rect 328454 539628 328460 539640
rect 245804 539600 328460 539628
rect 245804 539588 245810 539600
rect 328454 539588 328460 539600
rect 328512 539588 328518 539640
rect 245746 539452 245752 539504
rect 245804 539492 245810 539504
rect 245930 539492 245936 539504
rect 245804 539464 245936 539492
rect 245804 539452 245810 539464
rect 245930 539452 245936 539464
rect 245988 539452 245994 539504
rect 31570 538228 31576 538280
rect 31628 538268 31634 538280
rect 60734 538268 60740 538280
rect 31628 538240 60740 538268
rect 31628 538228 31634 538240
rect 60734 538228 60740 538240
rect 60792 538228 60798 538280
rect 257338 536800 257344 536852
rect 257396 536840 257402 536852
rect 579890 536840 579896 536852
rect 257396 536812 579896 536840
rect 257396 536800 257402 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 245838 536052 245844 536104
rect 245896 536092 245902 536104
rect 313274 536092 313280 536104
rect 245896 536064 313280 536092
rect 245896 536052 245902 536064
rect 313274 536052 313280 536064
rect 313332 536052 313338 536104
rect 57238 535440 57244 535492
rect 57296 535480 57302 535492
rect 60734 535480 60740 535492
rect 57296 535452 60740 535480
rect 57296 535440 57302 535452
rect 60734 535440 60740 535452
rect 60792 535440 60798 535492
rect 242986 532720 242992 532772
rect 243044 532760 243050 532772
rect 243262 532760 243268 532772
rect 243044 532732 243268 532760
rect 243044 532720 243050 532732
rect 243262 532720 243268 532732
rect 243320 532720 243326 532772
rect 46198 529864 46204 529916
rect 46256 529904 46262 529916
rect 53466 529904 53472 529916
rect 46256 529876 53472 529904
rect 46256 529864 46262 529876
rect 53466 529864 53472 529876
rect 53524 529864 53530 529916
rect 53466 528572 53472 528624
rect 53524 528612 53530 528624
rect 60734 528612 60740 528624
rect 53524 528584 60740 528612
rect 53524 528572 53530 528584
rect 60734 528572 60740 528584
rect 60792 528572 60798 528624
rect 3694 527144 3700 527196
rect 3752 527184 3758 527196
rect 4062 527184 4068 527196
rect 3752 527156 4068 527184
rect 3752 527144 3758 527156
rect 4062 527144 4068 527156
rect 4120 527184 4126 527196
rect 46198 527184 46204 527196
rect 4120 527156 46204 527184
rect 4120 527144 4126 527156
rect 46198 527144 46204 527156
rect 46256 527144 46262 527196
rect 245838 525784 245844 525836
rect 245896 525824 245902 525836
rect 282178 525824 282184 525836
rect 245896 525796 282184 525824
rect 245896 525784 245902 525796
rect 282178 525784 282184 525796
rect 282236 525784 282242 525836
rect 59170 521636 59176 521688
rect 59228 521676 59234 521688
rect 61654 521676 61660 521688
rect 59228 521648 61660 521676
rect 59228 521636 59234 521648
rect 61654 521636 61660 521648
rect 61712 521636 61718 521688
rect 245838 521636 245844 521688
rect 245896 521676 245902 521688
rect 349246 521676 349252 521688
rect 245896 521648 349252 521676
rect 245896 521636 245902 521648
rect 349246 521636 349252 521648
rect 349304 521636 349310 521688
rect 245838 518916 245844 518968
rect 245896 518956 245902 518968
rect 259546 518956 259552 518968
rect 245896 518928 259552 518956
rect 245896 518916 245902 518928
rect 259546 518916 259552 518928
rect 259604 518916 259610 518968
rect 3418 516060 3424 516112
rect 3476 516100 3482 516112
rect 58710 516100 58716 516112
rect 3476 516072 58716 516100
rect 3476 516060 3482 516072
rect 58710 516060 58716 516072
rect 58768 516060 58774 516112
rect 38562 514768 38568 514820
rect 38620 514808 38626 514820
rect 60734 514808 60740 514820
rect 38620 514780 60740 514808
rect 38620 514768 38626 514780
rect 60734 514768 60740 514780
rect 60792 514768 60798 514820
rect 245378 514768 245384 514820
rect 245436 514808 245442 514820
rect 263594 514808 263600 514820
rect 245436 514780 263600 514808
rect 245436 514768 245442 514780
rect 263594 514768 263600 514780
rect 263652 514768 263658 514820
rect 58710 513884 58716 513936
rect 58768 513924 58774 513936
rect 60090 513924 60096 513936
rect 58768 513896 60096 513924
rect 58768 513884 58774 513896
rect 60090 513884 60096 513896
rect 60148 513884 60154 513936
rect 245838 512592 245844 512644
rect 245896 512632 245902 512644
rect 251082 512632 251088 512644
rect 245896 512604 251088 512632
rect 245896 512592 245902 512604
rect 251082 512592 251088 512604
rect 251140 512632 251146 512644
rect 296714 512632 296720 512644
rect 251140 512604 296720 512632
rect 251140 512592 251146 512604
rect 296714 512592 296720 512604
rect 296772 512592 296778 512644
rect 251818 510620 251824 510672
rect 251876 510660 251882 510672
rect 580166 510660 580172 510672
rect 251876 510632 580172 510660
rect 251876 510620 251882 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 246666 509804 246672 509856
rect 246724 509844 246730 509856
rect 248322 509844 248328 509856
rect 246724 509816 248328 509844
rect 246724 509804 246730 509816
rect 248322 509804 248328 509816
rect 248380 509804 248386 509856
rect 248322 509260 248328 509312
rect 248380 509300 248386 509312
rect 249886 509300 249892 509312
rect 248380 509272 249892 509300
rect 248380 509260 248386 509272
rect 249886 509260 249892 509272
rect 249944 509260 249950 509312
rect 245838 506404 245844 506456
rect 245896 506444 245902 506456
rect 263686 506444 263692 506456
rect 245896 506416 263692 506444
rect 245896 506404 245902 506416
rect 263686 506404 263692 506416
rect 263744 506404 263750 506456
rect 263686 505724 263692 505776
rect 263744 505764 263750 505776
rect 300854 505764 300860 505776
rect 263744 505736 300860 505764
rect 263744 505724 263750 505736
rect 300854 505724 300860 505736
rect 300912 505724 300918 505776
rect 245838 502324 245844 502376
rect 245896 502364 245902 502376
rect 324958 502364 324964 502376
rect 245896 502336 324964 502364
rect 245896 502324 245902 502336
rect 324958 502324 324964 502336
rect 325016 502324 325022 502376
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 50430 501004 50436 501016
rect 3108 500976 50436 501004
rect 3108 500964 3114 500976
rect 50430 500964 50436 500976
rect 50488 500964 50494 501016
rect 55858 500964 55864 501016
rect 55916 501004 55922 501016
rect 60734 501004 60740 501016
rect 55916 500976 60740 501004
rect 55916 500964 55922 500976
rect 60734 500964 60740 500976
rect 60792 500964 60798 501016
rect 245838 499536 245844 499588
rect 245896 499576 245902 499588
rect 329834 499576 329840 499588
rect 245896 499548 329840 499576
rect 245896 499536 245902 499548
rect 329834 499536 329840 499548
rect 329892 499536 329898 499588
rect 262122 496816 262128 496868
rect 262180 496856 262186 496868
rect 304994 496856 305000 496868
rect 262180 496828 305000 496856
rect 262180 496816 262186 496828
rect 304994 496816 305000 496828
rect 305052 496816 305058 496868
rect 245838 496748 245844 496800
rect 245896 496788 245902 496800
rect 262140 496788 262168 496816
rect 245896 496760 262168 496788
rect 245896 496748 245902 496760
rect 48038 495456 48044 495508
rect 48096 495496 48102 495508
rect 60734 495496 60740 495508
rect 48096 495468 60740 495496
rect 48096 495456 48102 495468
rect 60734 495456 60740 495468
rect 60792 495456 60798 495508
rect 245838 492668 245844 492720
rect 245896 492708 245902 492720
rect 270494 492708 270500 492720
rect 245896 492680 270500 492708
rect 245896 492668 245902 492680
rect 270494 492668 270500 492680
rect 270552 492668 270558 492720
rect 56226 491308 56232 491360
rect 56284 491348 56290 491360
rect 60734 491348 60740 491360
rect 56284 491320 60740 491348
rect 56284 491308 56290 491320
rect 60734 491308 60740 491320
rect 60792 491308 60798 491360
rect 32950 488520 32956 488572
rect 33008 488560 33014 488572
rect 60734 488560 60740 488572
rect 33008 488532 60740 488560
rect 33008 488520 33014 488532
rect 60734 488520 60740 488532
rect 60792 488520 60798 488572
rect 43990 485800 43996 485852
rect 44048 485840 44054 485852
rect 61194 485840 61200 485852
rect 44048 485812 61200 485840
rect 44048 485800 44054 485812
rect 61194 485800 61200 485812
rect 61252 485800 61258 485852
rect 245838 485800 245844 485852
rect 245896 485840 245902 485852
rect 261478 485840 261484 485852
rect 245896 485812 261484 485840
rect 245896 485800 245902 485812
rect 261478 485800 261484 485812
rect 261536 485800 261542 485852
rect 251910 485732 251916 485784
rect 251968 485772 251974 485784
rect 580166 485772 580172 485784
rect 251968 485744 580172 485772
rect 251968 485732 251974 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 251082 482264 251088 482316
rect 251140 482304 251146 482316
rect 580258 482304 580264 482316
rect 251140 482276 580264 482304
rect 251140 482264 251146 482276
rect 580258 482264 580264 482276
rect 580316 482264 580322 482316
rect 59078 481652 59084 481704
rect 59136 481692 59142 481704
rect 61562 481692 61568 481704
rect 59136 481664 61568 481692
rect 59136 481652 59142 481664
rect 61562 481652 61568 481664
rect 61620 481652 61626 481704
rect 13078 477504 13084 477556
rect 13136 477544 13142 477556
rect 60734 477544 60740 477556
rect 13136 477516 60740 477544
rect 13136 477504 13142 477516
rect 60734 477504 60740 477516
rect 60792 477504 60798 477556
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 22738 474756 22744 474768
rect 3476 474728 22744 474756
rect 3476 474716 3482 474728
rect 22738 474716 22744 474728
rect 22796 474716 22802 474768
rect 245838 474716 245844 474768
rect 245896 474756 245902 474768
rect 317414 474756 317420 474768
rect 245896 474728 317420 474756
rect 245896 474716 245902 474728
rect 317414 474716 317420 474728
rect 317472 474716 317478 474768
rect 299474 472608 299480 472660
rect 299532 472648 299538 472660
rect 364334 472648 364340 472660
rect 299532 472620 364340 472648
rect 299532 472608 299538 472620
rect 364334 472608 364340 472620
rect 364392 472608 364398 472660
rect 245838 471996 245844 472048
rect 245896 472036 245902 472048
rect 299474 472036 299480 472048
rect 245896 472008 299480 472036
rect 245896 471996 245902 472008
rect 299474 471996 299480 472008
rect 299532 471996 299538 472048
rect 45370 470568 45376 470620
rect 45428 470608 45434 470620
rect 60918 470608 60924 470620
rect 45428 470580 60924 470608
rect 45428 470568 45434 470580
rect 60918 470568 60924 470580
rect 60976 470568 60982 470620
rect 275278 470568 275284 470620
rect 275336 470608 275342 470620
rect 580074 470608 580080 470620
rect 275336 470580 580080 470608
rect 275336 470568 275342 470580
rect 580074 470568 580080 470580
rect 580132 470568 580138 470620
rect 37090 467848 37096 467900
rect 37148 467888 37154 467900
rect 60734 467888 60740 467900
rect 37148 467860 60740 467888
rect 37148 467848 37154 467860
rect 60734 467848 60740 467860
rect 60792 467848 60798 467900
rect 53742 464992 53748 465044
rect 53800 465032 53806 465044
rect 60734 465032 60740 465044
rect 53800 465004 60740 465032
rect 53800 464992 53806 465004
rect 60734 464992 60740 465004
rect 60792 464992 60798 465044
rect 3418 463632 3424 463684
rect 3476 463672 3482 463684
rect 50338 463672 50344 463684
rect 3476 463644 50344 463672
rect 3476 463632 3482 463644
rect 50338 463632 50344 463644
rect 50396 463632 50402 463684
rect 17218 460912 17224 460964
rect 17276 460952 17282 460964
rect 52086 460952 52092 460964
rect 17276 460924 52092 460952
rect 17276 460912 17282 460924
rect 52086 460912 52092 460924
rect 52144 460952 52150 460964
rect 60734 460952 60740 460964
rect 52144 460924 60740 460952
rect 52144 460912 52150 460924
rect 60734 460912 60740 460924
rect 60792 460912 60798 460964
rect 245930 460912 245936 460964
rect 245988 460952 245994 460964
rect 269758 460952 269764 460964
rect 245988 460924 269764 460952
rect 245988 460912 245994 460924
rect 269758 460912 269764 460924
rect 269816 460912 269822 460964
rect 245930 458804 245936 458856
rect 245988 458844 245994 458856
rect 249978 458844 249984 458856
rect 245988 458816 249984 458844
rect 245988 458804 245994 458816
rect 249978 458804 249984 458816
rect 250036 458804 250042 458856
rect 50798 456764 50804 456816
rect 50856 456804 50862 456816
rect 60734 456804 60740 456816
rect 50856 456776 60740 456804
rect 50856 456764 50862 456776
rect 60734 456764 60740 456776
rect 60792 456764 60798 456816
rect 249058 456764 249064 456816
rect 249116 456804 249122 456816
rect 580166 456804 580172 456816
rect 249116 456776 580172 456804
rect 249116 456764 249122 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 245930 455404 245936 455456
rect 245988 455444 245994 455456
rect 263686 455444 263692 455456
rect 245988 455416 263692 455444
rect 245988 455404 245994 455416
rect 263686 455404 263692 455416
rect 263744 455404 263750 455456
rect 60642 455336 60648 455388
rect 60700 455376 60706 455388
rect 61378 455376 61384 455388
rect 60700 455348 61384 455376
rect 60700 455336 60706 455348
rect 61378 455336 61384 455348
rect 61436 455336 61442 455388
rect 246298 450508 246304 450560
rect 246356 450548 246362 450560
rect 252646 450548 252652 450560
rect 246356 450520 252652 450548
rect 246356 450508 246362 450520
rect 252646 450508 252652 450520
rect 252704 450508 252710 450560
rect 63218 449896 63224 449948
rect 63276 449936 63282 449948
rect 63494 449936 63500 449948
rect 63276 449908 63500 449936
rect 63276 449896 63282 449908
rect 63494 449896 63500 449908
rect 63552 449896 63558 449948
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 17218 449868 17224 449880
rect 3384 449840 17224 449868
rect 3384 449828 3390 449840
rect 17218 449828 17224 449840
rect 17276 449828 17282 449880
rect 245930 448536 245936 448588
rect 245988 448576 245994 448588
rect 255406 448576 255412 448588
rect 245988 448548 255412 448576
rect 245988 448536 245994 448548
rect 255406 448536 255412 448548
rect 255464 448536 255470 448588
rect 245378 447040 245384 447092
rect 245436 447080 245442 447092
rect 278038 447080 278044 447092
rect 245436 447052 278044 447080
rect 245436 447040 245442 447052
rect 278038 447040 278044 447052
rect 278096 447040 278102 447092
rect 54846 444388 54852 444440
rect 54904 444428 54910 444440
rect 60734 444428 60740 444440
rect 54904 444400 60740 444428
rect 54904 444388 54910 444400
rect 60734 444388 60740 444400
rect 60792 444388 60798 444440
rect 50890 441600 50896 441652
rect 50948 441640 50954 441652
rect 60734 441640 60740 441652
rect 50948 441612 60740 441640
rect 50948 441600 50954 441612
rect 60734 441600 60740 441612
rect 60792 441600 60798 441652
rect 245930 438880 245936 438932
rect 245988 438920 245994 438932
rect 278038 438920 278044 438932
rect 245988 438892 278044 438920
rect 245988 438880 245994 438892
rect 278038 438880 278044 438892
rect 278096 438880 278102 438932
rect 46658 437452 46664 437504
rect 46716 437492 46722 437504
rect 60918 437492 60924 437504
rect 46716 437464 60924 437492
rect 46716 437452 46722 437464
rect 60918 437452 60924 437464
rect 60976 437452 60982 437504
rect 59262 434732 59268 434784
rect 59320 434772 59326 434784
rect 61562 434772 61568 434784
rect 59320 434744 61568 434772
rect 59320 434732 59326 434744
rect 61562 434732 61568 434744
rect 61620 434732 61626 434784
rect 245930 434732 245936 434784
rect 245988 434772 245994 434784
rect 327258 434772 327264 434784
rect 245988 434744 327264 434772
rect 245988 434732 245994 434744
rect 327258 434732 327264 434744
rect 327316 434732 327322 434784
rect 251082 433344 251088 433356
rect 250824 433316 251088 433344
rect 57698 433236 57704 433288
rect 57756 433276 57762 433288
rect 62850 433276 62856 433288
rect 57756 433248 62856 433276
rect 57756 433236 57762 433248
rect 62850 433236 62856 433248
rect 62908 433236 62914 433288
rect 245930 433236 245936 433288
rect 245988 433276 245994 433288
rect 250824 433276 250852 433316
rect 251082 433304 251088 433316
rect 251140 433344 251146 433356
rect 306374 433344 306380 433356
rect 251140 433316 306380 433344
rect 251140 433304 251146 433316
rect 306374 433304 306380 433316
rect 306432 433304 306438 433356
rect 245988 433248 250852 433276
rect 245988 433236 245994 433248
rect 22738 428408 22744 428460
rect 22796 428448 22802 428460
rect 49418 428448 49424 428460
rect 22796 428420 49424 428448
rect 22796 428408 22802 428420
rect 49418 428408 49424 428420
rect 49476 428408 49482 428460
rect 49418 427796 49424 427848
rect 49476 427836 49482 427848
rect 60734 427836 60740 427848
rect 49476 427808 60740 427836
rect 49476 427796 49482 427808
rect 60734 427796 60740 427808
rect 60792 427796 60798 427848
rect 245930 427796 245936 427848
rect 245988 427836 245994 427848
rect 291930 427836 291936 427848
rect 245988 427808 291936 427836
rect 245988 427796 245994 427808
rect 291930 427796 291936 427808
rect 291988 427796 291994 427848
rect 252462 425688 252468 425740
rect 252520 425728 252526 425740
rect 291838 425728 291844 425740
rect 252520 425700 291844 425728
rect 252520 425688 252526 425700
rect 291838 425688 291844 425700
rect 291896 425688 291902 425740
rect 245930 425076 245936 425128
rect 245988 425116 245994 425128
rect 251358 425116 251364 425128
rect 245988 425088 251364 425116
rect 245988 425076 245994 425088
rect 251358 425076 251364 425088
rect 251416 425116 251422 425128
rect 252462 425116 252468 425128
rect 251416 425088 252468 425116
rect 251416 425076 251422 425088
rect 252462 425076 252468 425088
rect 252520 425076 252526 425128
rect 39758 423648 39764 423700
rect 39816 423688 39822 423700
rect 60734 423688 60740 423700
rect 39816 423660 60740 423688
rect 39816 423648 39822 423660
rect 60734 423648 60740 423660
rect 60792 423648 60798 423700
rect 245930 420928 245936 420980
rect 245988 420968 245994 420980
rect 322934 420968 322940 420980
rect 245988 420940 322940 420968
rect 245988 420928 245994 420940
rect 322934 420928 322940 420940
rect 322992 420928 322998 420980
rect 500218 419432 500224 419484
rect 500276 419472 500282 419484
rect 580166 419472 580172 419484
rect 500276 419444 580172 419472
rect 500276 419432 500282 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 245930 418208 245936 418260
rect 245988 418248 245994 418260
rect 247310 418248 247316 418260
rect 245988 418220 247316 418248
rect 245988 418208 245994 418220
rect 247310 418208 247316 418220
rect 247368 418208 247374 418260
rect 58986 417392 58992 417444
rect 59044 417432 59050 417444
rect 59998 417432 60004 417444
rect 59044 417404 60004 417432
rect 59044 417392 59050 417404
rect 59998 417392 60004 417404
rect 60056 417392 60062 417444
rect 62850 417392 62856 417444
rect 62908 417432 62914 417444
rect 63126 417432 63132 417444
rect 62908 417404 63132 417432
rect 62908 417392 62914 417404
rect 63126 417392 63132 417404
rect 63184 417392 63190 417444
rect 17218 416780 17224 416832
rect 17276 416820 17282 416832
rect 62298 416820 62304 416832
rect 17276 416792 62304 416820
rect 17276 416780 17282 416792
rect 62298 416780 62304 416792
rect 62356 416820 62362 416832
rect 63218 416820 63224 416832
rect 62356 416792 63224 416820
rect 62356 416780 62362 416792
rect 63218 416780 63224 416792
rect 63276 416780 63282 416832
rect 60458 416712 60464 416764
rect 60516 416752 60522 416764
rect 62758 416752 62764 416764
rect 60516 416724 62764 416752
rect 60516 416712 60522 416724
rect 62758 416712 62764 416724
rect 62816 416712 62822 416764
rect 42518 413992 42524 414044
rect 42576 414032 42582 414044
rect 60734 414032 60740 414044
rect 42576 414004 60740 414032
rect 42576 413992 42582 414004
rect 60734 413992 60740 414004
rect 60792 413992 60798 414044
rect 245930 413992 245936 414044
rect 245988 414032 245994 414044
rect 292758 414032 292764 414044
rect 245988 414004 292764 414032
rect 245988 413992 245994 414004
rect 292758 413992 292764 414004
rect 292816 413992 292822 414044
rect 245930 411272 245936 411324
rect 245988 411312 245994 411324
rect 298186 411312 298192 411324
rect 245988 411284 298192 411312
rect 245988 411272 245994 411284
rect 298186 411272 298192 411284
rect 298244 411272 298250 411324
rect 3418 411204 3424 411256
rect 3476 411244 3482 411256
rect 48958 411244 48964 411256
rect 3476 411216 48964 411244
rect 3476 411204 3482 411216
rect 48958 411204 48964 411216
rect 49016 411204 49022 411256
rect 53558 409980 53564 410032
rect 53616 410020 53622 410032
rect 53742 410020 53748 410032
rect 53616 409992 53748 410020
rect 53616 409980 53622 409992
rect 53742 409980 53748 409992
rect 53800 409980 53806 410032
rect 245286 408484 245292 408536
rect 245344 408524 245350 408536
rect 310606 408524 310612 408536
rect 245344 408496 310612 408524
rect 245344 408484 245350 408496
rect 310606 408484 310612 408496
rect 310664 408484 310670 408536
rect 37182 407736 37188 407788
rect 37240 407776 37246 407788
rect 60734 407776 60740 407788
rect 37240 407748 60740 407776
rect 37240 407736 37246 407748
rect 60734 407736 60740 407748
rect 60792 407736 60798 407788
rect 249150 407736 249156 407788
rect 249208 407776 249214 407788
rect 580350 407776 580356 407788
rect 249208 407748 580356 407776
rect 249208 407736 249214 407748
rect 580350 407736 580356 407748
rect 580408 407736 580414 407788
rect 243078 407124 243084 407176
rect 243136 407164 243142 407176
rect 245654 407164 245660 407176
rect 243136 407136 245660 407164
rect 243136 407124 243142 407136
rect 245654 407124 245660 407136
rect 245712 407124 245718 407176
rect 3510 407056 3516 407108
rect 3568 407096 3574 407108
rect 7834 407096 7840 407108
rect 3568 407068 7840 407096
rect 3568 407056 3574 407068
rect 7834 407056 7840 407068
rect 7892 407056 7898 407108
rect 7834 405696 7840 405748
rect 7892 405736 7898 405748
rect 8202 405736 8208 405748
rect 7892 405708 8208 405736
rect 7892 405696 7898 405708
rect 8202 405696 8208 405708
rect 8260 405736 8266 405748
rect 57330 405736 57336 405748
rect 8260 405708 57336 405736
rect 8260 405696 8266 405708
rect 57330 405696 57336 405708
rect 57388 405696 57394 405748
rect 53742 405084 53748 405136
rect 53800 405124 53806 405136
rect 66898 405124 66904 405136
rect 53800 405096 66904 405124
rect 53800 405084 53806 405096
rect 66898 405084 66904 405096
rect 66956 405084 66962 405136
rect 236638 405084 236644 405136
rect 236696 405124 236702 405136
rect 260834 405124 260840 405136
rect 236696 405096 260840 405124
rect 236696 405084 236702 405096
rect 260834 405084 260840 405096
rect 260892 405084 260898 405136
rect 56410 405016 56416 405068
rect 56468 405056 56474 405068
rect 80054 405056 80060 405068
rect 56468 405028 80060 405056
rect 56468 405016 56474 405028
rect 80054 405016 80060 405028
rect 80112 405016 80118 405068
rect 171042 405016 171048 405068
rect 171100 405056 171106 405068
rect 243078 405056 243084 405068
rect 171100 405028 243084 405056
rect 171100 405016 171106 405028
rect 243078 405016 243084 405028
rect 243136 405016 243142 405068
rect 57698 404948 57704 405000
rect 57756 404988 57762 405000
rect 104158 404988 104164 405000
rect 57756 404960 104164 404988
rect 57756 404948 57762 404960
rect 104158 404948 104164 404960
rect 104216 404948 104222 405000
rect 165522 404948 165528 405000
rect 165580 404988 165586 405000
rect 249886 404988 249892 405000
rect 165580 404960 249892 404988
rect 165580 404948 165586 404960
rect 249886 404948 249892 404960
rect 249944 404948 249950 405000
rect 8938 404472 8944 404524
rect 8996 404512 9002 404524
rect 96522 404512 96528 404524
rect 8996 404484 96528 404512
rect 8996 404472 9002 404484
rect 96522 404472 96528 404484
rect 96580 404512 96586 404524
rect 120718 404512 120724 404524
rect 96580 404484 120724 404512
rect 96580 404472 96586 404484
rect 120718 404472 120724 404484
rect 120776 404472 120782 404524
rect 202874 404472 202880 404524
rect 202932 404512 202938 404524
rect 203794 404512 203800 404524
rect 202932 404484 203800 404512
rect 202932 404472 202938 404484
rect 203794 404472 203800 404484
rect 203852 404512 203858 404524
rect 251818 404512 251824 404524
rect 203852 404484 251824 404512
rect 203852 404472 203858 404484
rect 251818 404472 251824 404484
rect 251876 404472 251882 404524
rect 50430 404404 50436 404456
rect 50488 404444 50494 404456
rect 178034 404444 178040 404456
rect 50488 404416 178040 404444
rect 50488 404404 50494 404416
rect 178034 404404 178040 404416
rect 178092 404404 178098 404456
rect 197354 404404 197360 404456
rect 197412 404444 197418 404456
rect 249058 404444 249064 404456
rect 197412 404416 249064 404444
rect 197412 404404 197418 404416
rect 249058 404404 249064 404416
rect 249116 404404 249122 404456
rect 66162 404336 66168 404388
rect 66220 404376 66226 404388
rect 580166 404376 580172 404388
rect 66220 404348 580172 404376
rect 66220 404336 66226 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 105262 404268 105268 404320
rect 105320 404308 105326 404320
rect 445018 404308 445024 404320
rect 105320 404280 445024 404308
rect 105320 404268 105326 404280
rect 445018 404268 445024 404280
rect 445076 404268 445082 404320
rect 14458 404200 14464 404252
rect 14516 404240 14522 404252
rect 242158 404240 242164 404252
rect 14516 404212 242164 404240
rect 14516 404200 14522 404212
rect 242158 404200 242164 404212
rect 242216 404200 242222 404252
rect 222838 404132 222844 404184
rect 222896 404172 222902 404184
rect 257338 404172 257344 404184
rect 222896 404144 257344 404172
rect 222896 404132 222902 404144
rect 257338 404132 257344 404144
rect 257396 404132 257402 404184
rect 63494 403996 63500 404048
rect 63552 404036 63558 404048
rect 63954 404036 63960 404048
rect 63552 404008 63960 404036
rect 63552 403996 63558 404008
rect 63954 403996 63960 404008
rect 64012 403996 64018 404048
rect 50982 403792 50988 403844
rect 51040 403832 51046 403844
rect 68278 403832 68284 403844
rect 51040 403804 68284 403832
rect 51040 403792 51046 403804
rect 68278 403792 68284 403804
rect 68336 403792 68342 403844
rect 55030 403724 55036 403776
rect 55088 403764 55094 403776
rect 73798 403764 73804 403776
rect 55088 403736 73804 403764
rect 55088 403724 55094 403736
rect 73798 403724 73804 403736
rect 73856 403724 73862 403776
rect 60366 403656 60372 403708
rect 60424 403696 60430 403708
rect 98730 403696 98736 403708
rect 60424 403668 98736 403696
rect 60424 403656 60430 403668
rect 98730 403656 98736 403668
rect 98788 403656 98794 403708
rect 239398 403656 239404 403708
rect 239456 403696 239462 403708
rect 248414 403696 248420 403708
rect 239456 403668 248420 403696
rect 239456 403656 239462 403668
rect 248414 403656 248420 403668
rect 248472 403656 248478 403708
rect 63126 403588 63132 403640
rect 63184 403628 63190 403640
rect 124214 403628 124220 403640
rect 63184 403600 124220 403628
rect 63184 403588 63190 403600
rect 124214 403588 124220 403600
rect 124272 403588 124278 403640
rect 148410 403588 148416 403640
rect 148468 403628 148474 403640
rect 251266 403628 251272 403640
rect 148468 403600 251272 403628
rect 148468 403588 148474 403600
rect 251266 403588 251272 403600
rect 251324 403588 251330 403640
rect 240134 403520 240140 403572
rect 240192 403560 240198 403572
rect 244458 403560 244464 403572
rect 240192 403532 244464 403560
rect 240192 403520 240198 403532
rect 244458 403520 244464 403532
rect 244516 403520 244522 403572
rect 46198 402908 46204 402960
rect 46256 402948 46262 402960
rect 200758 402948 200764 402960
rect 46256 402920 200764 402948
rect 46256 402908 46262 402920
rect 200758 402908 200764 402920
rect 200816 402908 200822 402960
rect 209590 402908 209596 402960
rect 209648 402948 209654 402960
rect 256602 402948 256608 402960
rect 209648 402920 256608 402948
rect 209648 402908 209654 402920
rect 256602 402908 256608 402920
rect 256660 402908 256666 402960
rect 57330 402840 57336 402892
rect 57388 402880 57394 402892
rect 181438 402880 181444 402892
rect 57388 402852 181444 402880
rect 57388 402840 57394 402852
rect 181438 402840 181444 402852
rect 181496 402840 181502 402892
rect 43438 402772 43444 402824
rect 43496 402812 43502 402824
rect 79318 402812 79324 402824
rect 43496 402784 79324 402812
rect 43496 402772 43502 402784
rect 79318 402772 79324 402784
rect 79376 402772 79382 402824
rect 161934 402772 161940 402824
rect 161992 402812 161998 402824
rect 162762 402812 162768 402824
rect 161992 402784 162768 402812
rect 161992 402772 161998 402784
rect 162762 402772 162768 402784
rect 162820 402812 162826 402824
rect 249150 402812 249156 402824
rect 162820 402784 249156 402812
rect 162820 402772 162826 402784
rect 249150 402772 249156 402784
rect 249208 402772 249214 402824
rect 100662 402296 100668 402348
rect 100720 402336 100726 402348
rect 108482 402336 108488 402348
rect 100720 402308 108488 402336
rect 100720 402296 100726 402308
rect 108482 402296 108488 402308
rect 108540 402296 108546 402348
rect 117498 402296 117504 402348
rect 117556 402336 117562 402348
rect 126974 402336 126980 402348
rect 117556 402308 126980 402336
rect 117556 402296 117562 402308
rect 126974 402296 126980 402308
rect 127032 402296 127038 402348
rect 164142 402296 164148 402348
rect 164200 402336 164206 402348
rect 171594 402336 171600 402348
rect 164200 402308 171600 402336
rect 164200 402296 164206 402308
rect 171594 402296 171600 402308
rect 171652 402296 171658 402348
rect 193858 402296 193864 402348
rect 193916 402336 193922 402348
rect 252646 402336 252652 402348
rect 193916 402308 252652 402336
rect 193916 402296 193922 402308
rect 252646 402296 252652 402308
rect 252704 402296 252710 402348
rect 256602 402296 256608 402348
rect 256660 402336 256666 402348
rect 299566 402336 299572 402348
rect 256660 402308 299572 402336
rect 256660 402296 256666 402308
rect 299566 402296 299572 402308
rect 299624 402296 299630 402348
rect 102042 402228 102048 402280
rect 102100 402268 102106 402280
rect 122098 402268 122104 402280
rect 102100 402240 122104 402268
rect 102100 402228 102106 402240
rect 122098 402228 122104 402240
rect 122156 402228 122162 402280
rect 136818 402228 136824 402280
rect 136876 402268 136882 402280
rect 146294 402268 146300 402280
rect 136876 402240 146300 402268
rect 136876 402228 136882 402240
rect 146294 402228 146300 402240
rect 146352 402228 146358 402280
rect 168282 402228 168288 402280
rect 168340 402268 168346 402280
rect 197354 402268 197360 402280
rect 168340 402240 197360 402268
rect 168340 402228 168346 402240
rect 197354 402228 197360 402240
rect 197412 402228 197418 402280
rect 232130 402228 232136 402280
rect 232188 402268 232194 402280
rect 309134 402268 309140 402280
rect 232188 402240 309140 402268
rect 232188 402228 232194 402240
rect 309134 402228 309140 402240
rect 309192 402228 309198 402280
rect 102778 401752 102784 401804
rect 102836 401792 102842 401804
rect 105262 401792 105268 401804
rect 102836 401764 105268 401792
rect 102836 401752 102842 401764
rect 105262 401752 105268 401764
rect 105320 401752 105326 401804
rect 116578 401616 116584 401668
rect 116636 401656 116642 401668
rect 123938 401656 123944 401668
rect 116636 401628 123944 401656
rect 116636 401616 116642 401628
rect 123938 401616 123944 401628
rect 123996 401616 124002 401668
rect 127158 401616 127164 401668
rect 127216 401656 127222 401668
rect 128998 401656 129004 401668
rect 127216 401628 129004 401656
rect 127216 401616 127222 401628
rect 128998 401616 129004 401628
rect 129056 401616 129062 401668
rect 158070 401616 158076 401668
rect 158128 401656 158134 401668
rect 158714 401656 158720 401668
rect 158128 401628 158720 401656
rect 158128 401616 158134 401628
rect 158714 401616 158720 401628
rect 158772 401616 158778 401668
rect 214558 401004 214564 401056
rect 214616 401044 214622 401056
rect 247310 401044 247316 401056
rect 214616 401016 247316 401044
rect 214616 401004 214622 401016
rect 247310 401004 247316 401016
rect 247368 401004 247374 401056
rect 177850 400936 177856 400988
rect 177908 400976 177914 400988
rect 242986 400976 242992 400988
rect 177908 400948 242992 400976
rect 177908 400936 177914 400948
rect 242986 400936 242992 400948
rect 243044 400936 243050 400988
rect 48130 400868 48136 400920
rect 48188 400908 48194 400920
rect 82078 400908 82084 400920
rect 48188 400880 82084 400908
rect 48188 400868 48194 400880
rect 82078 400868 82084 400880
rect 82136 400868 82142 400920
rect 173710 400868 173716 400920
rect 173768 400908 173774 400920
rect 255314 400908 255320 400920
rect 173768 400880 255320 400908
rect 173768 400868 173774 400880
rect 255314 400868 255320 400880
rect 255372 400868 255378 400920
rect 82722 400120 82728 400172
rect 82780 400160 82786 400172
rect 477494 400160 477500 400172
rect 82780 400132 477500 400160
rect 82780 400120 82786 400132
rect 477494 400120 477500 400132
rect 477552 400120 477558 400172
rect 53558 400052 53564 400104
rect 53616 400092 53622 400104
rect 296806 400092 296812 400104
rect 53616 400064 296812 400092
rect 53616 400052 53622 400064
rect 296806 400052 296812 400064
rect 296864 400092 296870 400104
rect 297358 400092 297364 400104
rect 296864 400064 297364 400092
rect 296864 400052 296870 400064
rect 297358 400052 297364 400064
rect 297416 400052 297422 400104
rect 173802 399576 173808 399628
rect 173860 399616 173866 399628
rect 187694 399616 187700 399628
rect 173860 399588 187700 399616
rect 173860 399576 173866 399588
rect 187694 399576 187700 399588
rect 187752 399576 187758 399628
rect 52270 399508 52276 399560
rect 52328 399548 52334 399560
rect 84838 399548 84844 399560
rect 52328 399520 84844 399548
rect 52328 399508 52334 399520
rect 84838 399508 84844 399520
rect 84896 399508 84902 399560
rect 111058 399508 111064 399560
rect 111116 399548 111122 399560
rect 136634 399548 136640 399560
rect 111116 399520 136640 399548
rect 111116 399508 111122 399520
rect 136634 399508 136640 399520
rect 136692 399508 136698 399560
rect 156598 399508 156604 399560
rect 156656 399548 156662 399560
rect 174814 399548 174820 399560
rect 156656 399520 174820 399548
rect 156656 399508 156662 399520
rect 174814 399508 174820 399520
rect 174872 399508 174878 399560
rect 179782 399508 179788 399560
rect 179840 399548 179846 399560
rect 206370 399548 206376 399560
rect 179840 399520 206376 399548
rect 179840 399508 179846 399520
rect 206370 399508 206376 399520
rect 206428 399508 206434 399560
rect 61746 399440 61752 399492
rect 61804 399480 61810 399492
rect 120718 399480 120724 399492
rect 61804 399452 120724 399480
rect 61804 399440 61810 399452
rect 120718 399440 120724 399452
rect 120776 399440 120782 399492
rect 145558 399440 145564 399492
rect 145616 399480 145622 399492
rect 259546 399480 259552 399492
rect 145616 399452 259552 399480
rect 145616 399440 145622 399452
rect 259546 399440 259552 399452
rect 259604 399440 259610 399492
rect 95142 398760 95148 398812
rect 95200 398800 95206 398812
rect 96522 398800 96528 398812
rect 95200 398772 96528 398800
rect 95200 398760 95206 398772
rect 96522 398760 96528 398772
rect 96580 398760 96586 398812
rect 123478 398148 123484 398200
rect 123536 398188 123542 398200
rect 194134 398188 194140 398200
rect 123536 398160 194140 398188
rect 123536 398148 123542 398160
rect 194134 398148 194140 398160
rect 194192 398148 194198 398200
rect 194594 398148 194600 398200
rect 194652 398188 194658 398200
rect 256694 398188 256700 398200
rect 194652 398160 256700 398188
rect 194652 398148 194658 398160
rect 256694 398148 256700 398160
rect 256752 398148 256758 398200
rect 3970 398080 3976 398132
rect 4028 398120 4034 398132
rect 5442 398120 5448 398132
rect 4028 398092 5448 398120
rect 4028 398080 4034 398092
rect 5442 398080 5448 398092
rect 5500 398120 5506 398132
rect 25498 398120 25504 398132
rect 5500 398092 25504 398120
rect 5500 398080 5506 398092
rect 25498 398080 25504 398092
rect 25556 398080 25562 398132
rect 170950 398080 170956 398132
rect 171008 398120 171014 398132
rect 251358 398120 251364 398132
rect 171008 398092 251364 398120
rect 171008 398080 171014 398092
rect 251358 398080 251364 398092
rect 251416 398080 251422 398132
rect 39666 396924 39672 396976
rect 39724 396964 39730 396976
rect 64138 396964 64144 396976
rect 39724 396936 64144 396964
rect 39724 396924 39730 396936
rect 64138 396924 64144 396936
rect 64196 396924 64202 396976
rect 135898 396924 135904 396976
rect 135956 396964 135962 396976
rect 168374 396964 168380 396976
rect 135956 396936 168380 396964
rect 135956 396924 135962 396936
rect 168374 396924 168380 396936
rect 168432 396924 168438 396976
rect 45278 396856 45284 396908
rect 45336 396896 45342 396908
rect 75178 396896 75184 396908
rect 45336 396868 75184 396896
rect 45336 396856 45342 396868
rect 75178 396856 75184 396868
rect 75236 396856 75242 396908
rect 153102 396856 153108 396908
rect 153160 396896 153166 396908
rect 190914 396896 190920 396908
rect 153160 396868 190920 396896
rect 153160 396856 153166 396868
rect 190914 396856 190920 396868
rect 190972 396856 190978 396908
rect 63218 396788 63224 396840
rect 63276 396828 63282 396840
rect 98638 396828 98644 396840
rect 63276 396800 98644 396828
rect 63276 396788 63282 396800
rect 98638 396788 98644 396800
rect 98696 396788 98702 396840
rect 157978 396788 157984 396840
rect 158036 396828 158042 396840
rect 240134 396828 240140 396840
rect 158036 396800 240140 396828
rect 158036 396788 158042 396800
rect 240134 396788 240140 396800
rect 240192 396788 240198 396840
rect 59078 396720 59084 396772
rect 59136 396760 59142 396772
rect 140774 396760 140780 396772
rect 59136 396732 140780 396760
rect 59136 396720 59142 396732
rect 140774 396720 140780 396732
rect 140832 396760 140838 396772
rect 582374 396760 582380 396772
rect 140832 396732 582380 396760
rect 140832 396720 140838 396732
rect 582374 396720 582380 396732
rect 582432 396720 582438 396772
rect 202138 395428 202144 395480
rect 202196 395468 202202 395480
rect 247218 395468 247224 395480
rect 202196 395440 247224 395468
rect 202196 395428 202202 395440
rect 247218 395428 247224 395440
rect 247276 395428 247282 395480
rect 175182 395360 175188 395412
rect 175240 395400 175246 395412
rect 249794 395400 249800 395412
rect 175240 395372 249800 395400
rect 175240 395360 175246 395372
rect 249794 395360 249800 395372
rect 249852 395360 249858 395412
rect 52178 395292 52184 395344
rect 52236 395332 52242 395344
rect 86218 395332 86224 395344
rect 52236 395304 86224 395332
rect 52236 395292 52242 395304
rect 86218 395292 86224 395304
rect 86276 395292 86282 395344
rect 148318 395292 148324 395344
rect 148376 395332 148382 395344
rect 245838 395332 245844 395344
rect 148376 395304 245844 395332
rect 148376 395292 148382 395304
rect 245838 395292 245844 395304
rect 245896 395332 245902 395344
rect 319438 395332 319444 395344
rect 245896 395304 319444 395332
rect 245896 395292 245902 395304
rect 319438 395292 319444 395304
rect 319496 395292 319502 395344
rect 45278 394000 45284 394052
rect 45336 394040 45342 394052
rect 85574 394040 85580 394052
rect 45336 394012 85580 394040
rect 45336 394000 45342 394012
rect 85574 394000 85580 394012
rect 85632 394000 85638 394052
rect 181438 394000 181444 394052
rect 181496 394040 181502 394052
rect 241514 394040 241520 394052
rect 181496 394012 241520 394040
rect 181496 394000 181502 394012
rect 241514 394000 241520 394012
rect 241572 394000 241578 394052
rect 48130 393932 48136 393984
rect 48188 393972 48194 393984
rect 95234 393972 95240 393984
rect 48188 393944 95240 393972
rect 48188 393932 48194 393944
rect 95234 393932 95240 393944
rect 95292 393932 95298 393984
rect 124858 393932 124864 393984
rect 124916 393972 124922 393984
rect 224954 393972 224960 393984
rect 124916 393944 224960 393972
rect 124916 393932 124922 393944
rect 224954 393932 224960 393944
rect 225012 393932 225018 393984
rect 246298 393320 246304 393372
rect 246356 393360 246362 393372
rect 315298 393360 315304 393372
rect 246356 393332 315304 393360
rect 246356 393320 246362 393332
rect 315298 393320 315304 393332
rect 315356 393320 315362 393372
rect 166258 392640 166264 392692
rect 166316 392680 166322 392692
rect 246298 392680 246304 392692
rect 166316 392652 246304 392680
rect 166316 392640 166322 392652
rect 246298 392640 246304 392652
rect 246356 392640 246362 392692
rect 176470 392572 176476 392624
rect 176528 392612 176534 392624
rect 258074 392612 258080 392624
rect 176528 392584 258080 392612
rect 176528 392572 176534 392584
rect 258074 392572 258080 392584
rect 258132 392572 258138 392624
rect 149698 391960 149704 392012
rect 149756 392000 149762 392012
rect 212534 392000 212540 392012
rect 149756 391972 212540 392000
rect 149756 391960 149762 391972
rect 212534 391960 212540 391972
rect 212592 391960 212598 392012
rect 246390 391960 246396 392012
rect 246448 392000 246454 392012
rect 353294 392000 353300 392012
rect 246448 391972 353300 392000
rect 246448 391960 246454 391972
rect 353294 391960 353300 391972
rect 353352 391960 353358 392012
rect 44082 391280 44088 391332
rect 44140 391320 44146 391332
rect 88334 391320 88340 391332
rect 44140 391292 88340 391320
rect 44140 391280 44146 391292
rect 88334 391280 88340 391292
rect 88392 391280 88398 391332
rect 212534 391280 212540 391332
rect 212592 391320 212598 391332
rect 256694 391320 256700 391332
rect 212592 391292 256700 391320
rect 212592 391280 212598 391292
rect 256694 391280 256700 391292
rect 256752 391280 256758 391332
rect 52362 391212 52368 391264
rect 52420 391252 52426 391264
rect 97994 391252 98000 391264
rect 52420 391224 98000 391252
rect 52420 391212 52426 391224
rect 97994 391212 98000 391224
rect 98052 391212 98058 391264
rect 153838 391212 153844 391264
rect 153896 391252 153902 391264
rect 246390 391252 246396 391264
rect 153896 391224 246396 391252
rect 153896 391212 153902 391224
rect 246390 391212 246396 391224
rect 246448 391212 246454 391264
rect 41138 388424 41144 388476
rect 41196 388464 41202 388476
rect 75914 388464 75920 388476
rect 41196 388436 75920 388464
rect 41196 388424 41202 388436
rect 75914 388424 75920 388436
rect 75972 388424 75978 388476
rect 178034 388288 178040 388340
rect 178092 388328 178098 388340
rect 178678 388328 178684 388340
rect 178092 388300 178684 388328
rect 178092 388288 178098 388300
rect 178678 388288 178684 388300
rect 178736 388288 178742 388340
rect 162118 388220 162124 388272
rect 162176 388260 162182 388272
rect 162762 388260 162768 388272
rect 162176 388232 162768 388260
rect 162176 388220 162182 388232
rect 162762 388220 162768 388232
rect 162820 388220 162826 388272
rect 135990 387880 135996 387932
rect 136048 387920 136054 387932
rect 178034 387920 178040 387932
rect 136048 387892 178040 387920
rect 136048 387880 136054 387892
rect 178034 387880 178040 387892
rect 178092 387880 178098 387932
rect 162762 387812 162768 387864
rect 162820 387852 162826 387864
rect 293954 387852 293960 387864
rect 162820 387824 293960 387852
rect 162820 387812 162826 387824
rect 293954 387812 293960 387824
rect 294012 387812 294018 387864
rect 45462 387744 45468 387796
rect 45520 387784 45526 387796
rect 113174 387784 113180 387796
rect 45520 387756 113180 387784
rect 45520 387744 45526 387756
rect 113174 387744 113180 387756
rect 113232 387784 113238 387796
rect 114462 387784 114468 387796
rect 113232 387756 114468 387784
rect 113232 387744 113238 387756
rect 114462 387744 114468 387756
rect 114520 387744 114526 387796
rect 114462 387064 114468 387116
rect 114520 387104 114526 387116
rect 293034 387104 293040 387116
rect 114520 387076 293040 387104
rect 114520 387064 114526 387076
rect 293034 387064 293040 387076
rect 293092 387064 293098 387116
rect 234614 385636 234620 385688
rect 234672 385676 234678 385688
rect 323026 385676 323032 385688
rect 234672 385648 323032 385676
rect 234672 385636 234678 385648
rect 323026 385636 323032 385648
rect 323084 385636 323090 385688
rect 242158 384344 242164 384396
rect 242216 384384 242222 384396
rect 262214 384384 262220 384396
rect 242216 384356 262220 384384
rect 242216 384344 242222 384356
rect 262214 384344 262220 384356
rect 262272 384344 262278 384396
rect 79318 384276 79324 384328
rect 79376 384316 79382 384328
rect 121454 384316 121460 384328
rect 79376 384288 121460 384316
rect 79376 384276 79382 384288
rect 121454 384276 121460 384288
rect 121512 384276 121518 384328
rect 132402 384276 132408 384328
rect 132460 384316 132466 384328
rect 245746 384316 245752 384328
rect 132460 384288 245752 384316
rect 132460 384276 132466 384288
rect 245746 384276 245752 384288
rect 245804 384276 245810 384328
rect 121454 383664 121460 383716
rect 121512 383704 121518 383716
rect 234614 383704 234620 383716
rect 121512 383676 234620 383704
rect 121512 383664 121518 383676
rect 234614 383664 234620 383676
rect 234672 383664 234678 383716
rect 63862 382916 63868 382968
rect 63920 382956 63926 382968
rect 138014 382956 138020 382968
rect 63920 382928 138020 382956
rect 63920 382916 63926 382928
rect 138014 382916 138020 382928
rect 138072 382916 138078 382968
rect 138014 382236 138020 382288
rect 138072 382276 138078 382288
rect 273898 382276 273904 382288
rect 138072 382248 273904 382276
rect 138072 382236 138078 382248
rect 273898 382236 273904 382248
rect 273956 382276 273962 382288
rect 275278 382276 275284 382288
rect 273956 382248 275284 382276
rect 273956 382236 273962 382248
rect 275278 382236 275284 382248
rect 275336 382236 275342 382288
rect 178678 381556 178684 381608
rect 178736 381596 178742 381608
rect 294046 381596 294052 381608
rect 178736 381568 294052 381596
rect 178736 381556 178742 381568
rect 294046 381556 294052 381568
rect 294104 381556 294110 381608
rect 126238 381488 126244 381540
rect 126296 381528 126302 381540
rect 255406 381528 255412 381540
rect 126296 381500 255412 381528
rect 126296 381488 126302 381500
rect 255406 381488 255412 381500
rect 255464 381488 255470 381540
rect 271322 379448 271328 379500
rect 271380 379488 271386 379500
rect 580166 379488 580172 379500
rect 271380 379460 580172 379488
rect 271380 379448 271386 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 217318 378768 217324 378820
rect 217376 378808 217382 378820
rect 270494 378808 270500 378820
rect 217376 378780 270500 378808
rect 217376 378768 217382 378780
rect 270494 378768 270500 378780
rect 270552 378808 270558 378820
rect 271322 378808 271328 378820
rect 270552 378780 271328 378808
rect 270552 378768 270558 378780
rect 271322 378768 271328 378780
rect 271380 378768 271386 378820
rect 218054 378088 218060 378140
rect 218112 378128 218118 378140
rect 251174 378128 251180 378140
rect 218112 378100 251180 378128
rect 218112 378088 218118 378100
rect 251174 378088 251180 378100
rect 251232 378128 251238 378140
rect 252462 378128 252468 378140
rect 251232 378100 252468 378128
rect 251232 378088 251238 378100
rect 252462 378088 252468 378100
rect 252520 378088 252526 378140
rect 60550 377408 60556 377460
rect 60608 377448 60614 377460
rect 109678 377448 109684 377460
rect 60608 377420 109684 377448
rect 60608 377408 60614 377420
rect 109678 377408 109684 377420
rect 109736 377408 109742 377460
rect 166810 377408 166816 377460
rect 166868 377448 166874 377460
rect 248506 377448 248512 377460
rect 166868 377420 248512 377448
rect 166868 377408 166874 377420
rect 248506 377408 248512 377420
rect 248564 377408 248570 377460
rect 252462 377408 252468 377460
rect 252520 377448 252526 377460
rect 270494 377448 270500 377460
rect 252520 377420 270500 377448
rect 252520 377408 252526 377420
rect 270494 377408 270500 377420
rect 270552 377408 270558 377460
rect 278038 377408 278044 377460
rect 278096 377448 278102 377460
rect 287054 377448 287060 377460
rect 278096 377420 287060 377448
rect 278096 377408 278102 377420
rect 287054 377408 287060 377420
rect 287112 377408 287118 377460
rect 220078 376048 220084 376100
rect 220136 376088 220142 376100
rect 247034 376088 247040 376100
rect 220136 376060 247040 376088
rect 220136 376048 220142 376060
rect 247034 376048 247040 376060
rect 247092 376048 247098 376100
rect 111702 375980 111708 376032
rect 111760 376020 111766 376032
rect 236638 376020 236644 376032
rect 111760 375992 236644 376020
rect 111760 375980 111766 375992
rect 236638 375980 236644 375992
rect 236696 375980 236702 376032
rect 91094 375300 91100 375352
rect 91152 375340 91158 375352
rect 92382 375340 92388 375352
rect 91152 375312 92388 375340
rect 91152 375300 91158 375312
rect 92382 375300 92388 375312
rect 92440 375300 92446 375352
rect 160830 374620 160836 374672
rect 160888 374660 160894 374672
rect 264974 374660 264980 374672
rect 160888 374632 264980 374660
rect 160888 374620 160894 374632
rect 264974 374620 264980 374632
rect 265032 374620 265038 374672
rect 92382 374008 92388 374060
rect 92440 374048 92446 374060
rect 295610 374048 295616 374060
rect 92440 374020 295616 374048
rect 92440 374008 92446 374020
rect 295610 374008 295616 374020
rect 295668 374008 295674 374060
rect 205634 373328 205640 373380
rect 205692 373368 205698 373380
rect 253198 373368 253204 373380
rect 205692 373340 253204 373368
rect 205692 373328 205698 373340
rect 253198 373328 253204 373340
rect 253256 373328 253262 373380
rect 59170 373260 59176 373312
rect 59228 373300 59234 373312
rect 113818 373300 113824 373312
rect 59228 373272 113824 373300
rect 59228 373260 59234 373272
rect 113818 373260 113824 373272
rect 113876 373260 113882 373312
rect 137278 373260 137284 373312
rect 137336 373300 137342 373312
rect 183554 373300 183560 373312
rect 137336 373272 183560 373300
rect 137336 373260 137342 373272
rect 183554 373260 183560 373272
rect 183612 373300 183618 373312
rect 231118 373300 231124 373312
rect 183612 373272 231124 373300
rect 183612 373260 183618 373272
rect 231118 373260 231124 373272
rect 231176 373260 231182 373312
rect 261478 373260 261484 373312
rect 261536 373300 261542 373312
rect 295518 373300 295524 373312
rect 261536 373272 295524 373300
rect 261536 373260 261542 373272
rect 295518 373260 295524 373272
rect 295576 373260 295582 373312
rect 164234 372580 164240 372632
rect 164292 372620 164298 372632
rect 164878 372620 164884 372632
rect 164292 372592 164884 372620
rect 164292 372580 164298 372592
rect 164878 372580 164884 372592
rect 164936 372620 164942 372632
rect 356054 372620 356060 372632
rect 164936 372592 356060 372620
rect 164936 372580 164942 372592
rect 356054 372580 356060 372592
rect 356112 372580 356118 372632
rect 43898 372172 43904 372224
rect 43956 372212 43962 372224
rect 44818 372212 44824 372224
rect 43956 372184 44824 372212
rect 43956 372172 43962 372184
rect 44818 372172 44824 372184
rect 44876 372172 44882 372224
rect 53650 371900 53656 371952
rect 53708 371940 53714 371952
rect 112438 371940 112444 371952
rect 53708 371912 112444 371940
rect 53708 371900 53714 371912
rect 112438 371900 112444 371912
rect 112496 371900 112502 371952
rect 209038 371900 209044 371952
rect 209096 371940 209102 371952
rect 217318 371940 217324 371952
rect 209096 371912 217324 371940
rect 209096 371900 209102 371912
rect 217318 371900 217324 371912
rect 217376 371900 217382 371952
rect 49418 371832 49424 371884
rect 49476 371872 49482 371884
rect 129826 371872 129832 371884
rect 49476 371844 129832 371872
rect 49476 371832 49482 371844
rect 129826 371832 129832 371844
rect 129884 371832 129890 371884
rect 215294 371832 215300 371884
rect 215352 371872 215358 371884
rect 279418 371872 279424 371884
rect 215352 371844 279424 371872
rect 215352 371832 215358 371844
rect 279418 371832 279424 371844
rect 279476 371832 279482 371884
rect 282178 371832 282184 371884
rect 282236 371872 282242 371884
rect 295334 371872 295340 371884
rect 282236 371844 295340 371872
rect 282236 371832 282242 371844
rect 295334 371832 295340 371844
rect 295392 371832 295398 371884
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 43898 371260 43904 371272
rect 3476 371232 43904 371260
rect 3476 371220 3482 371232
rect 43898 371220 43904 371232
rect 43956 371220 43962 371272
rect 129826 371220 129832 371272
rect 129884 371260 129890 371272
rect 202966 371260 202972 371272
rect 129884 371232 202972 371260
rect 129884 371220 129890 371232
rect 202966 371220 202972 371232
rect 203024 371220 203030 371272
rect 200758 370608 200764 370660
rect 200816 370648 200822 370660
rect 264974 370648 264980 370660
rect 200816 370620 264980 370648
rect 200816 370608 200822 370620
rect 264974 370608 264980 370620
rect 265032 370608 265038 370660
rect 168190 370540 168196 370592
rect 168248 370580 168254 370592
rect 239398 370580 239404 370592
rect 168248 370552 239404 370580
rect 168248 370540 168254 370552
rect 239398 370540 239404 370552
rect 239456 370540 239462 370592
rect 139302 370472 139308 370524
rect 139360 370512 139366 370524
rect 227714 370512 227720 370524
rect 139360 370484 227720 370512
rect 139360 370472 139366 370484
rect 227714 370472 227720 370484
rect 227772 370472 227778 370524
rect 243354 369180 243360 369232
rect 243412 369220 243418 369232
rect 252554 369220 252560 369232
rect 243412 369192 252560 369220
rect 243412 369180 243418 369192
rect 252554 369180 252560 369192
rect 252612 369180 252618 369232
rect 178678 369112 178684 369164
rect 178736 369152 178742 369164
rect 237374 369152 237380 369164
rect 178736 369124 237380 369152
rect 178736 369112 178742 369124
rect 237374 369112 237380 369124
rect 237432 369152 237438 369164
rect 294138 369152 294144 369164
rect 237432 369124 294144 369152
rect 237432 369112 237438 369124
rect 294138 369112 294144 369124
rect 294196 369112 294202 369164
rect 39666 368500 39672 368552
rect 39724 368540 39730 368552
rect 242986 368540 242992 368552
rect 39724 368512 242992 368540
rect 39724 368500 39730 368512
rect 242986 368500 242992 368512
rect 243044 368540 243050 368552
rect 243354 368540 243360 368552
rect 243044 368512 243360 368540
rect 243044 368500 243050 368512
rect 243354 368500 243360 368512
rect 243412 368500 243418 368552
rect 211798 367820 211804 367872
rect 211856 367860 211862 367872
rect 244550 367860 244556 367872
rect 211856 367832 244556 367860
rect 211856 367820 211862 367832
rect 244550 367820 244556 367832
rect 244608 367820 244614 367872
rect 129734 367752 129740 367804
rect 129792 367792 129798 367804
rect 143534 367792 143540 367804
rect 129792 367764 143540 367792
rect 129792 367752 129798 367764
rect 143534 367752 143540 367764
rect 143592 367792 143598 367804
rect 144270 367792 144276 367804
rect 143592 367764 144276 367792
rect 143592 367752 143598 367764
rect 144270 367752 144276 367764
rect 144328 367752 144334 367804
rect 169110 367752 169116 367804
rect 169168 367792 169174 367804
rect 263686 367792 263692 367804
rect 169168 367764 263692 367792
rect 169168 367752 169174 367764
rect 263686 367752 263692 367764
rect 263744 367752 263750 367804
rect 144270 367072 144276 367124
rect 144328 367112 144334 367124
rect 205634 367112 205640 367124
rect 144328 367084 205640 367112
rect 144328 367072 144334 367084
rect 205634 367072 205640 367084
rect 205692 367072 205698 367124
rect 52086 366392 52092 366444
rect 52144 366432 52150 366444
rect 70578 366432 70584 366444
rect 52144 366404 70584 366432
rect 52144 366392 52150 366404
rect 70578 366392 70584 366404
rect 70636 366392 70642 366444
rect 53466 366324 53472 366376
rect 53524 366364 53530 366376
rect 171962 366364 171968 366376
rect 53524 366336 171968 366364
rect 53524 366324 53530 366336
rect 171962 366324 171968 366336
rect 172020 366324 172026 366376
rect 152458 365780 152464 365832
rect 152516 365820 152522 365832
rect 276014 365820 276020 365832
rect 152516 365792 276020 365820
rect 152516 365780 152522 365792
rect 276014 365780 276020 365792
rect 276072 365780 276078 365832
rect 70578 365712 70584 365764
rect 70636 365752 70642 365764
rect 291286 365752 291292 365764
rect 70636 365724 291292 365752
rect 70636 365712 70642 365724
rect 291286 365712 291292 365724
rect 291344 365712 291350 365764
rect 54846 365032 54852 365084
rect 54904 365072 54910 365084
rect 96614 365072 96620 365084
rect 54904 365044 96620 365072
rect 54904 365032 54910 365044
rect 96614 365032 96620 365044
rect 96672 365032 96678 365084
rect 53742 364964 53748 365016
rect 53800 365004 53806 365016
rect 202874 365004 202880 365016
rect 53800 364976 202880 365004
rect 53800 364964 53806 364976
rect 202874 364964 202880 364976
rect 202932 365004 202938 365016
rect 301038 365004 301044 365016
rect 202932 364976 301044 365004
rect 202932 364964 202938 364976
rect 301038 364964 301044 364976
rect 301096 364964 301102 365016
rect 96614 364420 96620 364472
rect 96672 364460 96678 364472
rect 296898 364460 296904 364472
rect 96672 364432 296904 364460
rect 96672 364420 96678 364432
rect 296898 364420 296904 364432
rect 296956 364420 296962 364472
rect 158070 364352 158076 364404
rect 158128 364392 158134 364404
rect 160738 364392 160744 364404
rect 158128 364364 160744 364392
rect 158128 364352 158134 364364
rect 160738 364352 160744 364364
rect 160796 364352 160802 364404
rect 179230 364352 179236 364404
rect 179288 364392 179294 364404
rect 582374 364392 582380 364404
rect 179288 364364 582380 364392
rect 179288 364352 179294 364364
rect 582374 364352 582380 364364
rect 582432 364352 582438 364404
rect 160738 363740 160744 363792
rect 160796 363780 160802 363792
rect 245838 363780 245844 363792
rect 160796 363752 245844 363780
rect 160796 363740 160802 363752
rect 245838 363740 245844 363752
rect 245896 363740 245902 363792
rect 162210 363672 162216 363724
rect 162268 363712 162274 363724
rect 242802 363712 242808 363724
rect 162268 363684 242808 363712
rect 162268 363672 162274 363684
rect 242802 363672 242808 363684
rect 242860 363712 242866 363724
rect 347774 363712 347780 363724
rect 242860 363684 347780 363712
rect 242860 363672 242866 363684
rect 347774 363672 347780 363684
rect 347832 363672 347838 363724
rect 48038 363604 48044 363656
rect 48096 363644 48102 363656
rect 62114 363644 62120 363656
rect 48096 363616 62120 363644
rect 48096 363604 48102 363616
rect 62114 363604 62120 363616
rect 62172 363604 62178 363656
rect 144178 363604 144184 363656
rect 144236 363644 144242 363656
rect 178678 363644 178684 363656
rect 144236 363616 178684 363644
rect 144236 363604 144242 363616
rect 178678 363604 178684 363616
rect 178736 363604 178742 363656
rect 179322 363604 179328 363656
rect 179380 363644 179386 363656
rect 580902 363644 580908 363656
rect 179380 363616 580908 363644
rect 179380 363604 179386 363616
rect 580902 363604 580908 363616
rect 580960 363604 580966 363656
rect 62114 362924 62120 362976
rect 62172 362964 62178 362976
rect 62758 362964 62764 362976
rect 62172 362936 62764 362964
rect 62172 362924 62178 362936
rect 62758 362924 62764 362936
rect 62816 362964 62822 362976
rect 237466 362964 237472 362976
rect 62816 362936 237472 362964
rect 62816 362924 62822 362936
rect 237466 362924 237472 362936
rect 237524 362924 237530 362976
rect 240042 362924 240048 362976
rect 240100 362964 240106 362976
rect 310514 362964 310520 362976
rect 240100 362936 310520 362964
rect 240100 362924 240106 362936
rect 310514 362924 310520 362936
rect 310572 362924 310578 362976
rect 287698 362312 287704 362364
rect 287756 362352 287762 362364
rect 295426 362352 295432 362364
rect 287756 362324 295432 362352
rect 287756 362312 287762 362324
rect 295426 362312 295432 362324
rect 295484 362312 295490 362364
rect 55122 362176 55128 362228
rect 55180 362216 55186 362228
rect 100754 362216 100760 362228
rect 55180 362188 100760 362216
rect 55180 362176 55186 362188
rect 100754 362176 100760 362188
rect 100812 362176 100818 362228
rect 171778 361632 171784 361684
rect 171836 361672 171842 361684
rect 295518 361672 295524 361684
rect 171836 361644 295524 361672
rect 171836 361632 171842 361644
rect 295518 361632 295524 361644
rect 295576 361632 295582 361684
rect 100754 361564 100760 361616
rect 100812 361604 100818 361616
rect 298278 361604 298284 361616
rect 100812 361576 298284 361604
rect 100812 361564 100818 361576
rect 298278 361564 298284 361576
rect 298336 361564 298342 361616
rect 122742 360816 122748 360868
rect 122800 360856 122806 360868
rect 242894 360856 242900 360868
rect 122800 360828 242900 360856
rect 122800 360816 122806 360828
rect 242894 360816 242900 360828
rect 242952 360816 242958 360868
rect 250530 360408 250536 360460
rect 250588 360448 250594 360460
rect 309778 360448 309784 360460
rect 250588 360420 309784 360448
rect 250588 360408 250594 360420
rect 309778 360408 309784 360420
rect 309836 360408 309842 360460
rect 187418 360340 187424 360392
rect 187476 360380 187482 360392
rect 312538 360380 312544 360392
rect 187476 360352 312544 360380
rect 187476 360340 187482 360352
rect 312538 360340 312544 360352
rect 312596 360340 312602 360392
rect 31570 360272 31576 360324
rect 31628 360312 31634 360324
rect 302326 360312 302332 360324
rect 31628 360284 302332 360312
rect 31628 360272 31634 360284
rect 302326 360272 302332 360284
rect 302384 360272 302390 360324
rect 171870 360204 171876 360256
rect 171928 360244 171934 360256
rect 580258 360244 580264 360256
rect 171928 360216 580264 360244
rect 171928 360204 171934 360216
rect 580258 360204 580264 360216
rect 580316 360204 580322 360256
rect 163498 359456 163504 359508
rect 163556 359496 163562 359508
rect 193858 359496 193864 359508
rect 163556 359468 193864 359496
rect 163556 359456 163562 359468
rect 193858 359456 193864 359468
rect 193916 359456 193922 359508
rect 166902 358980 166908 359032
rect 166960 359020 166966 359032
rect 197722 359020 197728 359032
rect 166960 358992 197728 359020
rect 166960 358980 166966 358992
rect 197722 358980 197728 358992
rect 197780 358980 197786 359032
rect 172054 358912 172060 358964
rect 172112 358952 172118 358964
rect 220078 358952 220084 358964
rect 172112 358924 220084 358952
rect 172112 358912 172118 358924
rect 220078 358912 220084 358924
rect 220136 358952 220142 358964
rect 220262 358952 220268 358964
rect 220136 358924 220268 358952
rect 220136 358912 220142 358924
rect 220262 358912 220268 358924
rect 220320 358912 220326 358964
rect 129090 358844 129096 358896
rect 129148 358884 129154 358896
rect 202138 358884 202144 358896
rect 129148 358856 202144 358884
rect 129148 358844 129154 358856
rect 202138 358844 202144 358856
rect 202196 358844 202202 358896
rect 225414 358844 225420 358896
rect 225472 358884 225478 358896
rect 302234 358884 302240 358896
rect 225472 358856 302240 358884
rect 225472 358844 225478 358856
rect 302234 358844 302240 358856
rect 302292 358844 302298 358896
rect 181622 358776 181628 358828
rect 181680 358816 181686 358828
rect 337378 358816 337384 358828
rect 181680 358788 337384 358816
rect 181680 358776 181686 358788
rect 337378 358776 337384 358788
rect 337436 358776 337442 358828
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 17218 358748 17224 358760
rect 3384 358720 17224 358748
rect 3384 358708 3390 358720
rect 17218 358708 17224 358720
rect 17276 358708 17282 358760
rect 260098 358708 260104 358760
rect 260156 358748 260162 358760
rect 266630 358748 266636 358760
rect 260156 358720 266636 358748
rect 260156 358708 260162 358720
rect 266630 358708 266636 358720
rect 266688 358708 266694 358760
rect 290458 357756 290464 357808
rect 290516 357796 290522 357808
rect 308398 357796 308404 357808
rect 290516 357768 308404 357796
rect 290516 357756 290522 357768
rect 308398 357756 308404 357768
rect 308456 357756 308462 357808
rect 155862 357688 155868 357740
rect 155920 357728 155926 357740
rect 182910 357728 182916 357740
rect 155920 357700 182916 357728
rect 155920 357688 155926 357700
rect 182910 357688 182916 357700
rect 182968 357688 182974 357740
rect 282086 357688 282092 357740
rect 282144 357728 282150 357740
rect 313366 357728 313372 357740
rect 282144 357700 313372 357728
rect 282144 357688 282150 357700
rect 313366 357688 313372 357700
rect 313424 357688 313430 357740
rect 160002 357620 160008 357672
rect 160060 357660 160066 357672
rect 184934 357660 184940 357672
rect 160060 357632 184940 357660
rect 160060 357620 160066 357632
rect 184934 357620 184940 357632
rect 184992 357620 184998 357672
rect 260742 357620 260748 357672
rect 260800 357660 260806 357672
rect 305178 357660 305184 357672
rect 260800 357632 305184 357660
rect 260800 357620 260806 357632
rect 305178 357620 305184 357632
rect 305236 357620 305242 357672
rect 178770 357552 178776 357604
rect 178828 357592 178834 357604
rect 211798 357592 211804 357604
rect 178828 357564 211804 357592
rect 178828 357552 178834 357564
rect 211798 357552 211804 357564
rect 211856 357552 211862 357604
rect 223482 357552 223488 357604
rect 223540 357592 223546 357604
rect 298094 357592 298100 357604
rect 223540 357564 298100 357592
rect 223540 357552 223546 357564
rect 298094 357552 298100 357564
rect 298152 357552 298158 357604
rect 178678 357484 178684 357536
rect 178736 357524 178742 357536
rect 218330 357524 218336 357536
rect 178736 357496 218336 357524
rect 178736 357484 178742 357496
rect 218330 357484 218336 357496
rect 218388 357484 218394 357536
rect 227346 357484 227352 357536
rect 227404 357524 227410 357536
rect 342254 357524 342260 357536
rect 227404 357496 342260 357524
rect 227404 357484 227410 357496
rect 342254 357484 342260 357496
rect 342312 357484 342318 357536
rect 174630 357416 174636 357468
rect 174688 357456 174694 357468
rect 262214 357456 262220 357468
rect 174688 357428 262220 357456
rect 174688 357416 174694 357428
rect 262214 357416 262220 357428
rect 262272 357416 262278 357468
rect 279418 357416 279424 357468
rect 279476 357456 279482 357468
rect 449158 357456 449164 357468
rect 279476 357428 449164 357456
rect 279476 357416 279482 357428
rect 449158 357416 449164 357428
rect 449216 357416 449222 357468
rect 109034 357144 109040 357196
rect 109092 357184 109098 357196
rect 109678 357184 109684 357196
rect 109092 357156 109684 357184
rect 109092 357144 109098 357156
rect 109678 357144 109684 357156
rect 109736 357144 109742 357196
rect 193214 356776 193220 356788
rect 84166 356748 193220 356776
rect 55122 356668 55128 356720
rect 55180 356708 55186 356720
rect 80054 356708 80060 356720
rect 55180 356680 80060 356708
rect 55180 356668 55186 356680
rect 80054 356668 80060 356680
rect 80112 356708 80118 356720
rect 84166 356708 84194 356748
rect 193214 356736 193220 356748
rect 193272 356736 193278 356788
rect 80112 356680 84194 356708
rect 80112 356668 80118 356680
rect 109678 356668 109684 356720
rect 109736 356708 109742 356720
rect 254210 356708 254216 356720
rect 109736 356680 254216 356708
rect 109736 356668 109742 356680
rect 254210 356668 254216 356680
rect 254268 356668 254274 356720
rect 289078 356668 289084 356720
rect 289136 356708 289142 356720
rect 306466 356708 306472 356720
rect 289136 356680 306472 356708
rect 289136 356668 289142 356680
rect 306466 356668 306472 356680
rect 306524 356668 306530 356720
rect 171962 356260 171968 356312
rect 172020 356300 172026 356312
rect 199654 356300 199660 356312
rect 172020 356272 199660 356300
rect 172020 356260 172026 356272
rect 199654 356260 199660 356272
rect 199712 356260 199718 356312
rect 174538 356192 174544 356244
rect 174596 356232 174602 356244
rect 247126 356232 247132 356244
rect 174596 356204 247132 356232
rect 174596 356192 174602 356204
rect 247126 356192 247132 356204
rect 247184 356232 247190 356244
rect 247954 356232 247960 356244
rect 247184 356204 247960 356232
rect 247184 356192 247190 356204
rect 247954 356192 247960 356204
rect 248012 356192 248018 356244
rect 258902 356192 258908 356244
rect 258960 356232 258966 356244
rect 294230 356232 294236 356244
rect 258960 356204 294236 356232
rect 258960 356192 258966 356204
rect 294230 356192 294236 356204
rect 294288 356192 294294 356244
rect 117958 356124 117964 356176
rect 118016 356164 118022 356176
rect 214558 356164 214564 356176
rect 118016 356136 214564 356164
rect 118016 356124 118022 356136
rect 214558 356124 214564 356136
rect 214616 356124 214622 356176
rect 231118 356124 231124 356176
rect 231176 356164 231182 356176
rect 345658 356164 345664 356176
rect 231176 356136 345664 356164
rect 231176 356124 231182 356136
rect 345658 356124 345664 356136
rect 345716 356124 345722 356176
rect 46750 356056 46756 356108
rect 46808 356096 46814 356108
rect 305270 356096 305276 356108
rect 46808 356068 305276 356096
rect 46808 356056 46814 356068
rect 305270 356056 305276 356068
rect 305328 356056 305334 356108
rect 58986 355308 58992 355360
rect 59044 355348 59050 355360
rect 131114 355348 131120 355360
rect 59044 355320 131120 355348
rect 59044 355308 59050 355320
rect 131114 355308 131120 355320
rect 131172 355308 131178 355360
rect 194594 355240 194600 355292
rect 194652 355280 194658 355292
rect 195468 355280 195474 355292
rect 194652 355252 195474 355280
rect 194652 355240 194658 355252
rect 195468 355240 195474 355252
rect 195526 355240 195532 355292
rect 131114 355036 131120 355088
rect 131172 355076 131178 355088
rect 283374 355076 283380 355088
rect 131172 355048 283380 355076
rect 131172 355036 131178 355048
rect 283374 355036 283380 355048
rect 283432 355036 283438 355088
rect 165430 354968 165436 355020
rect 165488 355008 165494 355020
rect 209958 355008 209964 355020
rect 165488 354980 209964 355008
rect 165488 354968 165494 354980
rect 209958 354968 209964 354980
rect 210016 354968 210022 355020
rect 256970 354968 256976 355020
rect 257028 355008 257034 355020
rect 297358 355008 297364 355020
rect 257028 354980 297364 355008
rect 257028 354968 257034 354980
rect 297358 354968 297364 354980
rect 297416 354968 297422 355020
rect 179874 354900 179880 354952
rect 179932 354940 179938 354952
rect 287146 354940 287152 354952
rect 179932 354912 287152 354940
rect 179932 354900 179938 354912
rect 287146 354900 287152 354912
rect 287204 354940 287210 354952
rect 300118 354940 300124 354952
rect 287204 354912 300124 354940
rect 287204 354900 287210 354912
rect 300118 354900 300124 354912
rect 300176 354900 300182 354952
rect 170398 354832 170404 354884
rect 170456 354872 170462 354884
rect 279050 354872 279056 354884
rect 170456 354844 279056 354872
rect 170456 354832 170462 354844
rect 279050 354832 279056 354844
rect 279108 354832 279114 354884
rect 285950 354832 285956 354884
rect 286008 354872 286014 354884
rect 300946 354872 300952 354884
rect 286008 354844 300952 354872
rect 286008 354832 286014 354844
rect 300946 354832 300952 354844
rect 301004 354832 301010 354884
rect 68922 354764 68928 354816
rect 68980 354804 68986 354816
rect 194594 354804 194600 354816
rect 68980 354776 194600 354804
rect 68980 354764 68986 354776
rect 194594 354764 194600 354776
rect 194652 354764 194658 354816
rect 269022 354764 269028 354816
rect 269080 354804 269086 354816
rect 331490 354804 331496 354816
rect 269080 354776 331496 354804
rect 269080 354764 269086 354776
rect 331490 354764 331496 354776
rect 331548 354764 331554 354816
rect 275646 354696 275652 354748
rect 275704 354736 275710 354748
rect 305086 354736 305092 354748
rect 275704 354708 305092 354736
rect 275704 354696 275710 354708
rect 305086 354696 305092 354708
rect 305144 354696 305150 354748
rect 292298 354492 292304 354544
rect 292356 354532 292362 354544
rect 293310 354532 293316 354544
rect 292356 354504 293316 354532
rect 292356 354492 292362 354504
rect 293310 354492 293316 354504
rect 293368 354492 293374 354544
rect 175182 354356 175188 354408
rect 175240 354396 175246 354408
rect 176654 354396 176660 354408
rect 175240 354368 176660 354396
rect 175240 354356 175246 354368
rect 176654 354356 176660 354368
rect 176712 354356 176718 354408
rect 170858 352656 170864 352708
rect 170916 352696 170922 352708
rect 179782 352696 179788 352708
rect 170916 352668 179788 352696
rect 170916 352656 170922 352668
rect 179782 352656 179788 352668
rect 179840 352656 179846 352708
rect 90450 352588 90456 352640
rect 90508 352628 90514 352640
rect 178770 352628 178776 352640
rect 90508 352600 178776 352628
rect 90508 352588 90514 352600
rect 178770 352588 178776 352600
rect 178828 352588 178834 352640
rect 49418 352520 49424 352572
rect 49476 352560 49482 352572
rect 175182 352560 175188 352572
rect 49476 352532 175188 352560
rect 49476 352520 49482 352532
rect 175182 352520 175188 352532
rect 175240 352520 175246 352572
rect 175182 351908 175188 351960
rect 175240 351948 175246 351960
rect 177574 351948 177580 351960
rect 175240 351920 177580 351948
rect 175240 351908 175246 351920
rect 177574 351908 177580 351920
rect 177632 351908 177638 351960
rect 52086 351160 52092 351212
rect 52144 351200 52150 351212
rect 172054 351200 172060 351212
rect 52144 351172 172060 351200
rect 52144 351160 52150 351172
rect 172054 351160 172060 351172
rect 172112 351160 172118 351212
rect 50982 349800 50988 349852
rect 51040 349840 51046 349852
rect 152550 349840 152556 349852
rect 51040 349812 152556 349840
rect 51040 349800 51046 349812
rect 152550 349800 152556 349812
rect 152608 349800 152614 349852
rect 63402 348372 63408 348424
rect 63460 348412 63466 348424
rect 133966 348412 133972 348424
rect 63460 348384 133972 348412
rect 63460 348372 63466 348384
rect 133966 348372 133972 348384
rect 134024 348412 134030 348424
rect 134610 348412 134616 348424
rect 134024 348384 134616 348412
rect 134024 348372 134030 348384
rect 134610 348372 134616 348384
rect 134668 348372 134674 348424
rect 134610 347760 134616 347812
rect 134668 347800 134674 347812
rect 176654 347800 176660 347812
rect 134668 347772 176660 347800
rect 134668 347760 134674 347772
rect 176654 347760 176660 347772
rect 176712 347760 176718 347812
rect 14458 347012 14464 347064
rect 14516 347052 14522 347064
rect 35158 347052 35164 347064
rect 14516 347024 35164 347052
rect 14516 347012 14522 347024
rect 35158 347012 35164 347024
rect 35216 347012 35222 347064
rect 158622 345720 158628 345772
rect 158680 345760 158686 345772
rect 176654 345760 176660 345772
rect 158680 345732 176660 345760
rect 158680 345720 158686 345732
rect 176654 345720 176660 345732
rect 176712 345720 176718 345772
rect 3326 345652 3332 345704
rect 3384 345692 3390 345704
rect 14458 345692 14464 345704
rect 3384 345664 14464 345692
rect 3384 345652 3390 345664
rect 14458 345652 14464 345664
rect 14516 345652 14522 345704
rect 83458 345652 83464 345704
rect 83516 345692 83522 345704
rect 171778 345692 171784 345704
rect 83516 345664 171784 345692
rect 83516 345652 83522 345664
rect 171778 345652 171784 345664
rect 171836 345652 171842 345704
rect 295610 345652 295616 345704
rect 295668 345692 295674 345704
rect 468478 345692 468484 345704
rect 295668 345664 468484 345692
rect 295668 345652 295674 345664
rect 468478 345652 468484 345664
rect 468536 345652 468542 345704
rect 296070 343612 296076 343664
rect 296128 343652 296134 343664
rect 296714 343652 296720 343664
rect 296128 343624 296720 343652
rect 296128 343612 296134 343624
rect 296714 343612 296720 343624
rect 296772 343612 296778 343664
rect 126882 341504 126888 341556
rect 126940 341544 126946 341556
rect 179230 341544 179236 341556
rect 126940 341516 179236 341544
rect 126940 341504 126946 341516
rect 179230 341504 179236 341516
rect 179288 341544 179294 341556
rect 179506 341544 179512 341556
rect 179288 341516 179512 341544
rect 179288 341504 179294 341516
rect 179506 341504 179512 341516
rect 179564 341504 179570 341556
rect 132494 340892 132500 340944
rect 132552 340932 132558 340944
rect 132862 340932 132868 340944
rect 132552 340904 132868 340932
rect 132552 340892 132558 340904
rect 132862 340892 132868 340904
rect 132920 340932 132926 340944
rect 160738 340932 160744 340944
rect 132920 340904 160744 340932
rect 132920 340892 132926 340904
rect 160738 340892 160744 340904
rect 160796 340892 160802 340944
rect 75914 340144 75920 340196
rect 75972 340184 75978 340196
rect 132862 340184 132868 340196
rect 75972 340156 132868 340184
rect 75972 340144 75978 340156
rect 132862 340144 132868 340156
rect 132920 340144 132926 340196
rect 295610 339464 295616 339516
rect 295668 339504 295674 339516
rect 309870 339504 309876 339516
rect 295668 339476 309876 339504
rect 295668 339464 295674 339476
rect 309870 339464 309876 339476
rect 309928 339464 309934 339516
rect 295610 339124 295616 339176
rect 295668 339164 295674 339176
rect 298278 339164 298284 339176
rect 295668 339136 298284 339164
rect 295668 339124 295674 339136
rect 298278 339124 298284 339136
rect 298336 339124 298342 339176
rect 95050 338920 95056 338972
rect 95108 338960 95114 338972
rect 102778 338960 102784 338972
rect 95108 338932 102784 338960
rect 95108 338920 95114 338932
rect 102778 338920 102784 338932
rect 102836 338920 102842 338972
rect 163590 333956 163596 334008
rect 163648 333996 163654 334008
rect 176654 333996 176660 334008
rect 163648 333968 176660 333996
rect 163648 333956 163654 333968
rect 176654 333956 176660 333968
rect 176712 333956 176718 334008
rect 134518 333208 134524 333260
rect 134576 333248 134582 333260
rect 176470 333248 176476 333260
rect 134576 333220 176476 333248
rect 134576 333208 134582 333220
rect 176470 333208 176476 333220
rect 176528 333208 176534 333260
rect 157242 329808 157248 329860
rect 157300 329848 157306 329860
rect 176654 329848 176660 329860
rect 157300 329820 176660 329848
rect 157300 329808 157306 329820
rect 176654 329808 176660 329820
rect 176712 329808 176718 329860
rect 88334 329060 88340 329112
rect 88392 329100 88398 329112
rect 162210 329100 162216 329112
rect 88392 329072 162216 329100
rect 88392 329060 88398 329072
rect 162210 329060 162216 329072
rect 162268 329060 162274 329112
rect 295518 327700 295524 327752
rect 295576 327740 295582 327752
rect 347038 327740 347044 327752
rect 295576 327712 347044 327740
rect 295576 327700 295582 327712
rect 347038 327700 347044 327712
rect 347096 327700 347102 327752
rect 139486 327088 139492 327140
rect 139544 327128 139550 327140
rect 176654 327128 176660 327140
rect 139544 327100 176660 327128
rect 139544 327088 139550 327100
rect 176654 327088 176660 327100
rect 176712 327088 176718 327140
rect 325050 324300 325056 324352
rect 325108 324340 325114 324352
rect 580166 324340 580172 324352
rect 325108 324312 580172 324340
rect 325108 324300 325114 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 82722 323552 82728 323604
rect 82780 323592 82786 323604
rect 106274 323592 106280 323604
rect 82780 323564 106280 323592
rect 82780 323552 82786 323564
rect 106274 323552 106280 323564
rect 106332 323552 106338 323604
rect 66070 322192 66076 322244
rect 66128 322232 66134 322244
rect 164878 322232 164884 322244
rect 66128 322204 164884 322232
rect 66128 322192 66134 322204
rect 164878 322192 164884 322204
rect 164936 322192 164942 322244
rect 106274 321512 106280 321564
rect 106332 321552 106338 321564
rect 163590 321552 163596 321564
rect 106332 321524 163596 321552
rect 106332 321512 106338 321524
rect 163590 321512 163596 321524
rect 163648 321512 163654 321564
rect 295426 320152 295432 320204
rect 295484 320192 295490 320204
rect 335998 320192 336004 320204
rect 295484 320164 336004 320192
rect 295484 320152 295490 320164
rect 335998 320152 336004 320164
rect 336056 320152 336062 320204
rect 130470 319404 130476 319456
rect 130528 319444 130534 319456
rect 162118 319444 162124 319456
rect 130528 319416 162124 319444
rect 130528 319404 130534 319416
rect 162118 319404 162124 319416
rect 162176 319404 162182 319456
rect 3418 319064 3424 319116
rect 3476 319104 3482 319116
rect 8938 319104 8944 319116
rect 3476 319076 8944 319104
rect 3476 319064 3482 319076
rect 8938 319064 8944 319076
rect 8996 319064 9002 319116
rect 295426 318792 295432 318844
rect 295484 318832 295490 318844
rect 350534 318832 350540 318844
rect 295484 318804 350540 318832
rect 295484 318792 295490 318804
rect 350534 318792 350540 318804
rect 350592 318792 350598 318844
rect 100662 318112 100668 318164
rect 100720 318152 100726 318164
rect 133874 318152 133880 318164
rect 100720 318124 133880 318152
rect 100720 318112 100726 318124
rect 133874 318112 133880 318124
rect 133932 318112 133938 318164
rect 79318 318044 79324 318096
rect 79376 318084 79382 318096
rect 158070 318084 158076 318096
rect 79376 318056 158076 318084
rect 79376 318044 79382 318056
rect 158070 318044 158076 318056
rect 158128 318044 158134 318096
rect 295426 317364 295432 317416
rect 295484 317404 295490 317416
rect 302326 317404 302332 317416
rect 295484 317376 302332 317404
rect 295484 317364 295490 317376
rect 302326 317364 302332 317376
rect 302384 317364 302390 317416
rect 31570 316684 31576 316736
rect 31628 316724 31634 316736
rect 70486 316724 70492 316736
rect 31628 316696 70492 316724
rect 31628 316684 31634 316696
rect 70486 316684 70492 316696
rect 70544 316684 70550 316736
rect 302326 316684 302332 316736
rect 302384 316724 302390 316736
rect 467098 316724 467104 316736
rect 302384 316696 467104 316724
rect 302384 316684 302390 316696
rect 467098 316684 467104 316696
rect 467156 316684 467162 316736
rect 175090 316412 175096 316464
rect 175148 316452 175154 316464
rect 177574 316452 177580 316464
rect 175148 316424 177580 316452
rect 175148 316412 175154 316424
rect 177574 316412 177580 316424
rect 177632 316412 177638 316464
rect 169018 316044 169024 316056
rect 125566 316016 169024 316044
rect 73154 315936 73160 315988
rect 73212 315976 73218 315988
rect 125566 315976 125594 316016
rect 169018 316004 169024 316016
rect 169076 316004 169082 316056
rect 73212 315948 125594 315976
rect 73212 315936 73218 315948
rect 162762 315256 162768 315308
rect 162820 315296 162826 315308
rect 176654 315296 176660 315308
rect 162820 315268 176660 315296
rect 162820 315256 162826 315268
rect 176654 315256 176660 315268
rect 176712 315256 176718 315308
rect 71866 314644 71872 314696
rect 71924 314684 71930 314696
rect 73154 314684 73160 314696
rect 71924 314656 73160 314684
rect 71924 314644 71930 314656
rect 73154 314644 73160 314656
rect 73212 314644 73218 314696
rect 103606 314032 103612 314084
rect 103664 314072 103670 314084
rect 134518 314072 134524 314084
rect 103664 314044 134524 314072
rect 103664 314032 103670 314044
rect 134518 314032 134524 314044
rect 134576 314032 134582 314084
rect 49602 313964 49608 314016
rect 49660 314004 49666 314016
rect 126422 314004 126428 314016
rect 49660 313976 126428 314004
rect 49660 313964 49666 313976
rect 126422 313964 126428 313976
rect 126480 313964 126486 314016
rect 14458 313896 14464 313948
rect 14516 313936 14522 313948
rect 118694 313936 118700 313948
rect 14516 313908 118700 313936
rect 14516 313896 14522 313908
rect 118694 313896 118700 313908
rect 118752 313896 118758 313948
rect 293862 313284 293868 313336
rect 293920 313324 293926 313336
rect 356698 313324 356704 313336
rect 293920 313296 356704 313324
rect 293920 313284 293926 313296
rect 356698 313284 356704 313296
rect 356756 313284 356762 313336
rect 167730 313216 167736 313268
rect 167788 313256 167794 313268
rect 170950 313256 170956 313268
rect 167788 313228 170956 313256
rect 167788 313216 167794 313228
rect 170950 313216 170956 313228
rect 171008 313256 171014 313268
rect 176654 313256 176660 313268
rect 171008 313228 176660 313256
rect 171008 313216 171014 313228
rect 176654 313216 176660 313228
rect 176712 313216 176718 313268
rect 300118 313216 300124 313268
rect 300176 313256 300182 313268
rect 580166 313256 580172 313268
rect 300176 313228 580172 313256
rect 300176 313216 300182 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 8938 311788 8944 311840
rect 8996 311828 9002 311840
rect 41414 311828 41420 311840
rect 8996 311800 41420 311828
rect 8996 311788 9002 311800
rect 41414 311788 41420 311800
rect 41472 311788 41478 311840
rect 50798 311176 50804 311228
rect 50856 311216 50862 311228
rect 124306 311216 124312 311228
rect 50856 311188 124312 311216
rect 50856 311176 50862 311188
rect 124306 311176 124312 311188
rect 124364 311176 124370 311228
rect 41414 311108 41420 311160
rect 41472 311148 41478 311160
rect 42610 311148 42616 311160
rect 41472 311120 42616 311148
rect 41472 311108 41478 311120
rect 42610 311108 42616 311120
rect 42668 311148 42674 311160
rect 116670 311148 116676 311160
rect 42668 311120 116676 311148
rect 42668 311108 42674 311120
rect 116670 311108 116676 311120
rect 116728 311108 116734 311160
rect 295334 310428 295340 310480
rect 295392 310468 295398 310480
rect 305270 310468 305276 310480
rect 295392 310440 305276 310468
rect 295392 310428 295398 310440
rect 305270 310428 305276 310440
rect 305328 310468 305334 310480
rect 305454 310468 305460 310480
rect 305328 310440 305460 310468
rect 305328 310428 305334 310440
rect 305454 310428 305460 310440
rect 305512 310428 305518 310480
rect 116762 309816 116768 309868
rect 116820 309856 116826 309868
rect 176654 309856 176660 309868
rect 116820 309828 176660 309856
rect 116820 309816 116826 309828
rect 176654 309816 176660 309828
rect 176712 309816 176718 309868
rect 41230 309748 41236 309800
rect 41288 309788 41294 309800
rect 121546 309788 121552 309800
rect 41288 309760 121552 309788
rect 41288 309748 41294 309760
rect 121546 309748 121552 309760
rect 121604 309748 121610 309800
rect 305454 309748 305460 309800
rect 305512 309788 305518 309800
rect 355318 309788 355324 309800
rect 305512 309760 355324 309788
rect 305512 309748 305518 309760
rect 355318 309748 355324 309760
rect 355376 309748 355382 309800
rect 43990 308456 43996 308508
rect 44048 308496 44054 308508
rect 132494 308496 132500 308508
rect 44048 308468 132500 308496
rect 44048 308456 44054 308468
rect 132494 308456 132500 308468
rect 132552 308456 132558 308508
rect 33042 308388 33048 308440
rect 33100 308428 33106 308440
rect 127802 308428 127808 308440
rect 33100 308400 127808 308428
rect 33100 308388 33106 308400
rect 127802 308388 127808 308400
rect 127860 308388 127866 308440
rect 295518 308388 295524 308440
rect 295576 308428 295582 308440
rect 302326 308428 302332 308440
rect 295576 308400 302332 308428
rect 295576 308388 295582 308400
rect 302326 308388 302332 308400
rect 302384 308388 302390 308440
rect 97994 308116 98000 308168
rect 98052 308156 98058 308168
rect 98730 308156 98736 308168
rect 98052 308128 98736 308156
rect 98052 308116 98058 308128
rect 98730 308116 98736 308128
rect 98788 308116 98794 308168
rect 98730 307776 98736 307828
rect 98788 307816 98794 307828
rect 153930 307816 153936 307828
rect 98788 307788 153936 307816
rect 98788 307776 98794 307788
rect 153930 307776 153936 307788
rect 153988 307776 153994 307828
rect 81434 307368 81440 307420
rect 81492 307408 81498 307420
rect 82078 307408 82084 307420
rect 81492 307380 82084 307408
rect 81492 307368 81498 307380
rect 82078 307368 82084 307380
rect 82136 307368 82142 307420
rect 75178 306416 75184 306468
rect 75236 306456 75242 306468
rect 133138 306456 133144 306468
rect 75236 306428 133144 306456
rect 75236 306416 75242 306428
rect 133138 306416 133144 306428
rect 133196 306416 133202 306468
rect 81434 306348 81440 306400
rect 81492 306388 81498 306400
rect 142890 306388 142896 306400
rect 81492 306360 142896 306388
rect 81492 306348 81498 306360
rect 142890 306348 142896 306360
rect 142948 306348 142954 306400
rect 68278 305668 68284 305720
rect 68336 305708 68342 305720
rect 97258 305708 97264 305720
rect 68336 305680 97264 305708
rect 68336 305668 68342 305680
rect 97258 305668 97264 305680
rect 97316 305668 97322 305720
rect 46750 305600 46756 305652
rect 46808 305640 46814 305652
rect 80054 305640 80060 305652
rect 46808 305612 80060 305640
rect 46808 305600 46814 305612
rect 80054 305600 80060 305612
rect 80112 305600 80118 305652
rect 121362 305600 121368 305652
rect 121420 305640 121426 305652
rect 177850 305640 177856 305652
rect 121420 305612 177856 305640
rect 121420 305600 121426 305612
rect 177850 305600 177856 305612
rect 177908 305600 177914 305652
rect 86402 305056 86408 305108
rect 86460 305096 86466 305108
rect 131850 305096 131856 305108
rect 86460 305068 131856 305096
rect 86460 305056 86466 305068
rect 131850 305056 131856 305068
rect 131908 305056 131914 305108
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 120074 305028 120080 305040
rect 3292 305000 120080 305028
rect 3292 304988 3298 305000
rect 120074 304988 120080 305000
rect 120132 305028 120138 305040
rect 121362 305028 121368 305040
rect 120132 305000 121368 305028
rect 120132 304988 120138 305000
rect 121362 304988 121368 305000
rect 121420 304988 121426 305040
rect 68830 304240 68836 304292
rect 68888 304280 68894 304292
rect 174630 304280 174636 304292
rect 68888 304252 174636 304280
rect 68888 304240 68894 304252
rect 174630 304240 174636 304252
rect 174688 304240 174694 304292
rect 157150 303696 157156 303748
rect 157208 303736 157214 303748
rect 176654 303736 176660 303748
rect 157208 303708 176660 303736
rect 157208 303696 157214 303708
rect 176654 303696 176660 303708
rect 176712 303696 176718 303748
rect 114002 303628 114008 303680
rect 114060 303668 114066 303680
rect 171778 303668 171784 303680
rect 114060 303640 171784 303668
rect 114060 303628 114066 303640
rect 171778 303628 171784 303640
rect 171836 303628 171842 303680
rect 73798 303560 73804 303612
rect 73856 303600 73862 303612
rect 88978 303600 88984 303612
rect 73856 303572 88984 303600
rect 73856 303560 73862 303572
rect 88978 303560 88984 303572
rect 89036 303560 89042 303612
rect 111794 302948 111800 303000
rect 111852 302988 111858 303000
rect 132586 302988 132592 303000
rect 111852 302960 132592 302988
rect 111852 302948 111858 302960
rect 132586 302948 132592 302960
rect 132644 302948 132650 303000
rect 46842 302880 46848 302932
rect 46900 302920 46906 302932
rect 69474 302920 69480 302932
rect 46900 302892 69480 302920
rect 46900 302880 46906 302892
rect 69474 302880 69480 302892
rect 69532 302880 69538 302932
rect 92382 302880 92388 302932
rect 92440 302920 92446 302932
rect 115290 302920 115296 302932
rect 92440 302892 115296 302920
rect 92440 302880 92446 302892
rect 115290 302880 115296 302892
rect 115348 302880 115354 302932
rect 92842 302336 92848 302388
rect 92900 302376 92906 302388
rect 162118 302376 162124 302388
rect 92900 302348 162124 302376
rect 92900 302336 92906 302348
rect 162118 302336 162124 302348
rect 162176 302336 162182 302388
rect 59078 302268 59084 302320
rect 59136 302308 59142 302320
rect 145558 302308 145564 302320
rect 59136 302280 145564 302308
rect 59136 302268 59142 302280
rect 145558 302268 145564 302280
rect 145616 302308 145622 302320
rect 145742 302308 145748 302320
rect 145616 302280 145748 302308
rect 145616 302268 145622 302280
rect 145742 302268 145748 302280
rect 145800 302268 145806 302320
rect 69106 302200 69112 302252
rect 69164 302240 69170 302252
rect 69474 302240 69480 302252
rect 69164 302212 69480 302240
rect 69164 302200 69170 302212
rect 69474 302200 69480 302212
rect 69532 302240 69538 302252
rect 167638 302240 167644 302252
rect 69532 302212 167644 302240
rect 69532 302200 69538 302212
rect 167638 302200 167644 302212
rect 167696 302200 167702 302252
rect 110874 301520 110880 301572
rect 110932 301560 110938 301572
rect 111702 301560 111708 301572
rect 110932 301532 111708 301560
rect 110932 301520 110938 301532
rect 111702 301520 111708 301532
rect 111760 301560 111766 301572
rect 143626 301560 143632 301572
rect 111760 301532 143632 301560
rect 111760 301520 111766 301532
rect 143626 301520 143632 301532
rect 143684 301520 143690 301572
rect 91094 301452 91100 301504
rect 91152 301492 91158 301504
rect 167730 301492 167736 301504
rect 91152 301464 167736 301492
rect 91152 301452 91158 301464
rect 167730 301452 167736 301464
rect 167788 301452 167794 301504
rect 97258 300840 97264 300892
rect 97316 300880 97322 300892
rect 151078 300880 151084 300892
rect 97316 300852 151084 300880
rect 97316 300840 97322 300852
rect 151078 300840 151084 300852
rect 151136 300840 151142 300892
rect 295334 300840 295340 300892
rect 295392 300880 295398 300892
rect 305270 300880 305276 300892
rect 295392 300852 305276 300880
rect 295392 300840 295398 300852
rect 305270 300840 305276 300852
rect 305328 300840 305334 300892
rect 142154 300772 142160 300824
rect 142212 300812 142218 300824
rect 143442 300812 143448 300824
rect 142212 300784 143448 300812
rect 142212 300772 142218 300784
rect 143442 300772 143448 300784
rect 143500 300772 143506 300824
rect 94130 300568 94136 300620
rect 94188 300608 94194 300620
rect 95142 300608 95148 300620
rect 94188 300580 95148 300608
rect 94188 300568 94194 300580
rect 95142 300568 95148 300580
rect 95200 300568 95206 300620
rect 108298 299820 108304 299872
rect 108356 299860 108362 299872
rect 111794 299860 111800 299872
rect 108356 299832 111800 299860
rect 108356 299820 108362 299832
rect 111794 299820 111800 299832
rect 111852 299820 111858 299872
rect 84194 299752 84200 299804
rect 84252 299792 84258 299804
rect 142982 299792 142988 299804
rect 84252 299764 142988 299792
rect 84252 299752 84258 299764
rect 142982 299752 142988 299764
rect 143040 299752 143046 299804
rect 95142 299684 95148 299736
rect 95200 299724 95206 299736
rect 155310 299724 155316 299736
rect 95200 299696 155316 299724
rect 95200 299684 95206 299696
rect 155310 299684 155316 299696
rect 155368 299684 155374 299736
rect 79226 299616 79232 299668
rect 79284 299656 79290 299668
rect 159450 299656 159456 299668
rect 79284 299628 159456 299656
rect 79284 299616 79290 299628
rect 159450 299616 159456 299628
rect 159508 299616 159514 299668
rect 77386 299548 77392 299600
rect 77444 299588 77450 299600
rect 160830 299588 160836 299600
rect 77444 299560 160836 299588
rect 77444 299548 77450 299560
rect 160830 299548 160836 299560
rect 160888 299548 160894 299600
rect 32398 299480 32404 299532
rect 32456 299520 32462 299532
rect 117958 299520 117964 299532
rect 32456 299492 117964 299520
rect 32456 299480 32462 299492
rect 117958 299480 117964 299492
rect 118016 299480 118022 299532
rect 143442 299480 143448 299532
rect 143500 299520 143506 299532
rect 174630 299520 174636 299532
rect 143500 299492 174636 299520
rect 143500 299480 143506 299492
rect 174630 299480 174636 299492
rect 174688 299480 174694 299532
rect 166994 299412 167000 299464
rect 167052 299452 167058 299464
rect 168282 299452 168288 299464
rect 167052 299424 168288 299452
rect 167052 299412 167058 299424
rect 168282 299412 168288 299424
rect 168340 299452 168346 299464
rect 176654 299452 176660 299464
rect 168340 299424 176660 299452
rect 168340 299412 168346 299424
rect 176654 299412 176660 299424
rect 176712 299412 176718 299464
rect 297358 299412 297364 299464
rect 297416 299452 297422 299464
rect 580166 299452 580172 299464
rect 297416 299424 580172 299452
rect 297416 299412 297422 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 60458 298800 60464 298852
rect 60516 298840 60522 298852
rect 120166 298840 120172 298852
rect 60516 298812 120172 298840
rect 60516 298800 60522 298812
rect 120166 298800 120172 298812
rect 120224 298800 120230 298852
rect 53558 298732 53564 298784
rect 53616 298772 53622 298784
rect 166994 298772 167000 298784
rect 53616 298744 167000 298772
rect 53616 298732 53622 298744
rect 166994 298732 167000 298744
rect 167052 298732 167058 298784
rect 91738 298324 91744 298376
rect 91796 298364 91802 298376
rect 133230 298364 133236 298376
rect 91796 298336 133236 298364
rect 91796 298324 91802 298336
rect 133230 298324 133236 298336
rect 133288 298324 133294 298376
rect 106734 298256 106740 298308
rect 106792 298296 106798 298308
rect 148410 298296 148416 298308
rect 106792 298268 148416 298296
rect 106792 298256 106798 298268
rect 148410 298256 148416 298268
rect 148468 298256 148474 298308
rect 83550 298188 83556 298240
rect 83608 298228 83614 298240
rect 145558 298228 145564 298240
rect 83608 298200 145564 298228
rect 83608 298188 83614 298200
rect 145558 298188 145564 298200
rect 145616 298188 145622 298240
rect 66162 298120 66168 298172
rect 66220 298160 66226 298172
rect 140130 298160 140136 298172
rect 66220 298132 140136 298160
rect 66220 298120 66226 298132
rect 140130 298120 140136 298132
rect 140188 298120 140194 298172
rect 115934 298052 115940 298104
rect 115992 298092 115998 298104
rect 116578 298092 116584 298104
rect 115992 298064 116584 298092
rect 115992 298052 115998 298064
rect 116578 298052 116584 298064
rect 116636 298052 116642 298104
rect 8202 297440 8208 297492
rect 8260 297480 8266 297492
rect 72602 297480 72608 297492
rect 8260 297452 72608 297480
rect 8260 297440 8266 297452
rect 72602 297440 72608 297452
rect 72660 297440 72666 297492
rect 95050 297440 95056 297492
rect 95108 297480 95114 297492
rect 176654 297480 176660 297492
rect 95108 297452 176660 297480
rect 95108 297440 95114 297452
rect 176654 297440 176660 297452
rect 176712 297440 176718 297492
rect 43898 297372 43904 297424
rect 43956 297412 43962 297424
rect 129274 297412 129280 297424
rect 43956 297384 129280 297412
rect 43956 297372 43962 297384
rect 129274 297372 129280 297384
rect 129332 297372 129338 297424
rect 102226 296828 102232 296880
rect 102284 296868 102290 296880
rect 148502 296868 148508 296880
rect 102284 296840 148508 296868
rect 102284 296828 102290 296840
rect 148502 296828 148508 296840
rect 148560 296828 148566 296880
rect 90634 296760 90640 296812
rect 90692 296800 90698 296812
rect 138658 296800 138664 296812
rect 90692 296772 138664 296800
rect 90692 296760 90698 296772
rect 138658 296760 138664 296772
rect 138716 296760 138722 296812
rect 86126 296692 86132 296744
rect 86184 296732 86190 296744
rect 151170 296732 151176 296744
rect 86184 296704 151176 296732
rect 86184 296692 86190 296704
rect 151170 296692 151176 296704
rect 151228 296692 151234 296744
rect 115106 295672 115112 295724
rect 115164 295712 115170 295724
rect 116762 295712 116768 295724
rect 115164 295684 116768 295712
rect 115164 295672 115170 295684
rect 116762 295672 116768 295684
rect 116820 295672 116826 295724
rect 100938 295604 100944 295656
rect 100996 295644 101002 295656
rect 127618 295644 127624 295656
rect 100996 295616 127624 295644
rect 100996 295604 101002 295616
rect 127618 295604 127624 295616
rect 127676 295604 127682 295656
rect 88058 295536 88064 295588
rect 88116 295576 88122 295588
rect 126330 295576 126336 295588
rect 88116 295548 126336 295576
rect 88116 295536 88122 295548
rect 126330 295536 126336 295548
rect 126388 295536 126394 295588
rect 87414 295468 87420 295520
rect 87472 295508 87478 295520
rect 131758 295508 131764 295520
rect 87472 295480 131764 295508
rect 87472 295468 87478 295480
rect 131758 295468 131764 295480
rect 131816 295468 131822 295520
rect 43438 295400 43444 295452
rect 43496 295440 43502 295452
rect 100754 295440 100760 295452
rect 43496 295412 100760 295440
rect 43496 295400 43502 295412
rect 100754 295400 100760 295412
rect 100812 295440 100818 295452
rect 101582 295440 101588 295452
rect 100812 295412 101588 295440
rect 100812 295400 100818 295412
rect 101582 295400 101588 295412
rect 101640 295400 101646 295452
rect 110598 295400 110604 295452
rect 110656 295440 110662 295452
rect 149974 295440 149980 295452
rect 110656 295412 149980 295440
rect 110656 295400 110662 295412
rect 149974 295400 149980 295412
rect 150032 295400 150038 295452
rect 82262 295332 82268 295384
rect 82320 295372 82326 295384
rect 149790 295372 149796 295384
rect 82320 295344 149796 295372
rect 82320 295332 82326 295344
rect 149790 295332 149796 295344
rect 149848 295332 149854 295384
rect 295518 295332 295524 295384
rect 295576 295372 295582 295384
rect 300118 295372 300124 295384
rect 295576 295344 300124 295372
rect 295576 295332 295582 295344
rect 300118 295332 300124 295344
rect 300176 295332 300182 295384
rect 50890 295264 50896 295316
rect 50948 295304 50954 295316
rect 71774 295304 71780 295316
rect 50948 295276 71780 295304
rect 50948 295264 50954 295276
rect 71774 295264 71780 295276
rect 71832 295264 71838 295316
rect 174630 295264 174636 295316
rect 174688 295304 174694 295316
rect 176654 295304 176660 295316
rect 174688 295276 176660 295304
rect 174688 295264 174694 295276
rect 176654 295264 176660 295276
rect 176712 295264 176718 295316
rect 64138 294584 64144 294636
rect 64196 294624 64202 294636
rect 64690 294624 64696 294636
rect 64196 294596 64696 294624
rect 64196 294584 64202 294596
rect 64690 294584 64696 294596
rect 64748 294624 64754 294636
rect 70670 294624 70676 294636
rect 64748 294596 70676 294624
rect 64748 294584 64754 294596
rect 70670 294584 70676 294596
rect 70728 294584 70734 294636
rect 73246 294584 73252 294636
rect 73304 294624 73310 294636
rect 75178 294624 75184 294636
rect 73304 294596 75184 294624
rect 73304 294584 73310 294596
rect 75178 294584 75184 294596
rect 75236 294584 75242 294636
rect 95786 294584 95792 294636
rect 95844 294624 95850 294636
rect 173710 294624 173716 294636
rect 95844 294596 173716 294624
rect 95844 294584 95850 294596
rect 173710 294584 173716 294596
rect 173768 294584 173774 294636
rect 74534 294516 74540 294568
rect 74592 294556 74598 294568
rect 91738 294556 91744 294568
rect 74592 294528 91744 294556
rect 74592 294516 74598 294528
rect 91738 294516 91744 294528
rect 91796 294516 91802 294568
rect 89806 294176 89812 294228
rect 89864 294216 89870 294228
rect 95878 294216 95884 294228
rect 89864 294188 95884 294216
rect 89864 294176 89870 294188
rect 95878 294176 95884 294188
rect 95936 294216 95942 294228
rect 96430 294216 96436 294228
rect 95936 294188 96436 294216
rect 95936 294176 95942 294188
rect 96430 294176 96436 294188
rect 96488 294176 96494 294228
rect 105446 294176 105452 294228
rect 105504 294216 105510 294228
rect 115934 294216 115940 294228
rect 105504 294188 115940 294216
rect 105504 294176 105510 294188
rect 115934 294176 115940 294188
rect 115992 294216 115998 294228
rect 123662 294216 123668 294228
rect 115992 294188 123668 294216
rect 115992 294176 115998 294188
rect 123662 294176 123668 294188
rect 123720 294176 123726 294228
rect 59998 294108 60004 294160
rect 60056 294148 60062 294160
rect 92474 294148 92480 294160
rect 60056 294120 92480 294148
rect 60056 294108 60062 294120
rect 92474 294108 92480 294120
rect 92532 294108 92538 294160
rect 93854 294108 93860 294160
rect 93912 294148 93918 294160
rect 124950 294148 124956 294160
rect 93912 294120 124956 294148
rect 93912 294108 93918 294120
rect 124950 294108 124956 294120
rect 125008 294108 125014 294160
rect 79042 294080 79048 294092
rect 64846 294052 79048 294080
rect 4798 293972 4804 294024
rect 4856 294012 4862 294024
rect 64846 294012 64874 294052
rect 79042 294040 79048 294052
rect 79100 294080 79106 294092
rect 79318 294080 79324 294092
rect 79100 294052 79324 294080
rect 79100 294040 79106 294052
rect 79318 294040 79324 294052
rect 79376 294040 79382 294092
rect 80974 294040 80980 294092
rect 81032 294080 81038 294092
rect 117958 294080 117964 294092
rect 81032 294052 117964 294080
rect 81032 294040 81038 294052
rect 117958 294040 117964 294052
rect 118016 294040 118022 294092
rect 4856 293984 64874 294012
rect 4856 293972 4862 293984
rect 77110 293972 77116 294024
rect 77168 294012 77174 294024
rect 83458 294012 83464 294024
rect 77168 293984 83464 294012
rect 77168 293972 77174 293984
rect 83458 293972 83464 293984
rect 83516 293972 83522 294024
rect 85482 293972 85488 294024
rect 85540 294012 85546 294024
rect 90450 294012 90456 294024
rect 85540 293984 90456 294012
rect 85540 293972 85546 293984
rect 90450 293972 90456 293984
rect 90508 293972 90514 294024
rect 91922 293972 91928 294024
rect 91980 294012 91986 294024
rect 140038 294012 140044 294024
rect 91980 293984 140044 294012
rect 91980 293972 91986 293984
rect 140038 293972 140044 293984
rect 140096 293972 140102 294024
rect 295334 293972 295340 294024
rect 295392 294012 295398 294024
rect 307018 294012 307024 294024
rect 295392 293984 307024 294012
rect 295392 293972 295398 293984
rect 307018 293972 307024 293984
rect 307076 293972 307082 294024
rect 103606 293904 103612 293956
rect 103664 293944 103670 293956
rect 104526 293944 104532 293956
rect 103664 293916 104532 293944
rect 103664 293904 103670 293916
rect 104526 293904 104532 293916
rect 104584 293904 104590 293956
rect 109034 293904 109040 293956
rect 109092 293944 109098 293956
rect 109678 293944 109684 293956
rect 109092 293916 109684 293944
rect 109092 293904 109098 293916
rect 109678 293904 109684 293916
rect 109736 293904 109742 293956
rect 46842 293292 46848 293344
rect 46900 293332 46906 293344
rect 69014 293332 69020 293344
rect 46900 293304 69020 293332
rect 46900 293292 46906 293304
rect 69014 293292 69020 293304
rect 69072 293292 69078 293344
rect 2682 293224 2688 293276
rect 2740 293264 2746 293276
rect 89806 293264 89812 293276
rect 2740 293236 89812 293264
rect 2740 293224 2746 293236
rect 89806 293224 89812 293236
rect 89864 293224 89870 293276
rect 98362 293224 98368 293276
rect 98420 293264 98426 293276
rect 98638 293264 98644 293276
rect 98420 293236 98644 293264
rect 98420 293224 98426 293236
rect 98638 293224 98644 293236
rect 98696 293224 98702 293276
rect 68830 293088 68836 293140
rect 68888 293088 68894 293140
rect 68848 292936 68876 293088
rect 68830 292884 68836 292936
rect 68888 292884 68894 292936
rect 116670 292884 116676 292936
rect 116728 292924 116734 292936
rect 126514 292924 126520 292936
rect 116728 292896 126520 292924
rect 116728 292884 116734 292896
rect 126514 292884 126520 292896
rect 126572 292884 126578 292936
rect 92474 292816 92480 292868
rect 92532 292856 92538 292868
rect 123754 292856 123760 292868
rect 92532 292828 123760 292856
rect 92532 292816 92538 292828
rect 123754 292816 123760 292828
rect 123812 292816 123818 292868
rect 99650 292748 99656 292800
rect 99708 292788 99714 292800
rect 157978 292788 157984 292800
rect 99708 292760 157984 292788
rect 99708 292748 99714 292760
rect 157978 292748 157984 292760
rect 158036 292748 158042 292800
rect 75178 292680 75184 292732
rect 75236 292720 75242 292732
rect 136082 292720 136088 292732
rect 75236 292692 136088 292720
rect 75236 292680 75242 292692
rect 136082 292680 136088 292692
rect 136140 292680 136146 292732
rect 58618 292612 58624 292664
rect 58676 292652 58682 292664
rect 96706 292652 96712 292664
rect 58676 292624 96712 292652
rect 58676 292612 58682 292624
rect 96706 292612 96712 292624
rect 96764 292612 96770 292664
rect 98362 292612 98368 292664
rect 98420 292652 98426 292664
rect 174630 292652 174636 292664
rect 98420 292624 174636 292652
rect 98420 292612 98426 292624
rect 174630 292612 174636 292624
rect 174688 292612 174694 292664
rect 69198 292544 69204 292596
rect 69256 292584 69262 292596
rect 71958 292584 71964 292596
rect 69256 292556 71964 292584
rect 69256 292544 69262 292556
rect 71958 292544 71964 292556
rect 72016 292544 72022 292596
rect 84838 292544 84844 292596
rect 84896 292584 84902 292596
rect 176010 292584 176016 292596
rect 84896 292556 176016 292584
rect 84896 292544 84902 292556
rect 176010 292544 176016 292556
rect 176068 292544 176074 292596
rect 67450 291864 67456 291916
rect 67508 291904 67514 291916
rect 73706 291904 73712 291916
rect 67508 291876 73712 291904
rect 67508 291864 67514 291876
rect 73706 291864 73712 291876
rect 73764 291864 73770 291916
rect 83274 291864 83280 291916
rect 83332 291904 83338 291916
rect 83332 291876 84194 291904
rect 83332 291864 83338 291876
rect 2866 291388 2872 291440
rect 2924 291428 2930 291440
rect 8938 291428 8944 291440
rect 2924 291400 8944 291428
rect 2924 291388 2930 291400
rect 8938 291388 8944 291400
rect 8996 291388 9002 291440
rect 84166 291224 84194 291876
rect 103146 291864 103152 291916
rect 103204 291904 103210 291916
rect 103204 291876 103514 291904
rect 103204 291864 103210 291876
rect 103486 291292 103514 291876
rect 112806 291864 112812 291916
rect 112864 291904 112870 291916
rect 112864 291876 113174 291904
rect 112864 291864 112870 291876
rect 113146 291360 113174 291876
rect 117314 291864 117320 291916
rect 117372 291904 117378 291916
rect 120810 291904 120816 291916
rect 117372 291876 120816 291904
rect 117372 291864 117378 291876
rect 120810 291864 120816 291876
rect 120868 291864 120874 291916
rect 127710 291796 127716 291848
rect 127768 291836 127774 291848
rect 143442 291836 143448 291848
rect 127768 291808 143448 291836
rect 127768 291796 127774 291808
rect 143442 291796 143448 291808
rect 143500 291836 143506 291848
rect 163590 291836 163596 291848
rect 143500 291808 163596 291836
rect 143500 291796 143506 291808
rect 163590 291796 163596 291808
rect 163648 291796 163654 291848
rect 137370 291360 137376 291372
rect 113146 291332 137376 291360
rect 137370 291320 137376 291332
rect 137428 291320 137434 291372
rect 134610 291292 134616 291304
rect 103486 291264 134616 291292
rect 134610 291252 134616 291264
rect 134668 291252 134674 291304
rect 129182 291224 129188 291236
rect 84166 291196 129188 291224
rect 129182 291184 129188 291196
rect 129240 291184 129246 291236
rect 295610 291184 295616 291236
rect 295668 291224 295674 291236
rect 301222 291224 301228 291236
rect 295668 291196 301228 291224
rect 295668 291184 295674 291196
rect 301222 291184 301228 291196
rect 301280 291184 301286 291236
rect 166994 291116 167000 291168
rect 167052 291156 167058 291168
rect 168190 291156 168196 291168
rect 167052 291128 168196 291156
rect 167052 291116 167058 291128
rect 168190 291116 168196 291128
rect 168248 291156 168254 291168
rect 176654 291156 176660 291168
rect 168248 291128 176660 291156
rect 168248 291116 168254 291128
rect 176654 291116 176660 291128
rect 176712 291116 176718 291168
rect 295518 291116 295524 291168
rect 295576 291156 295582 291168
rect 301038 291156 301044 291168
rect 295576 291128 301044 291156
rect 295576 291116 295582 291128
rect 301038 291116 301044 291128
rect 301096 291116 301102 291168
rect 17218 290436 17224 290488
rect 17276 290476 17282 290488
rect 35802 290476 35808 290488
rect 17276 290448 35808 290476
rect 17276 290436 17282 290448
rect 35802 290436 35808 290448
rect 35860 290476 35866 290488
rect 52454 290476 52460 290488
rect 35860 290448 52460 290476
rect 35860 290436 35866 290448
rect 52454 290436 52460 290448
rect 52512 290436 52518 290488
rect 121454 289960 121460 290012
rect 121512 290000 121518 290012
rect 144270 290000 144276 290012
rect 121512 289972 144276 290000
rect 121512 289960 121518 289972
rect 144270 289960 144276 289972
rect 144328 289960 144334 290012
rect 52454 289892 52460 289944
rect 52512 289932 52518 289944
rect 53650 289932 53656 289944
rect 52512 289904 53656 289932
rect 52512 289892 52518 289904
rect 53650 289892 53656 289904
rect 53708 289932 53714 289944
rect 67726 289932 67732 289944
rect 53708 289904 67732 289932
rect 53708 289892 53714 289904
rect 67726 289892 67732 289904
rect 67784 289892 67790 289944
rect 121638 289892 121644 289944
rect 121696 289932 121702 289944
rect 149882 289932 149888 289944
rect 121696 289904 149888 289932
rect 121696 289892 121702 289904
rect 149882 289892 149888 289904
rect 149940 289892 149946 289944
rect 48038 289824 48044 289876
rect 48096 289864 48102 289876
rect 67634 289864 67640 289876
rect 48096 289836 67640 289864
rect 48096 289824 48102 289836
rect 67634 289824 67640 289836
rect 67692 289824 67698 289876
rect 172146 289864 172152 289876
rect 126900 289836 172152 289864
rect 121454 289756 121460 289808
rect 121512 289796 121518 289808
rect 126422 289796 126428 289808
rect 121512 289768 126428 289796
rect 121512 289756 121518 289768
rect 126422 289756 126428 289768
rect 126480 289796 126486 289808
rect 126900 289796 126928 289836
rect 172146 289824 172152 289836
rect 172204 289824 172210 289876
rect 126480 289768 126928 289796
rect 126480 289756 126486 289768
rect 35802 289076 35808 289128
rect 35860 289116 35866 289128
rect 67726 289116 67732 289128
rect 35860 289088 67732 289116
rect 35860 289076 35866 289088
rect 67726 289076 67732 289088
rect 67784 289076 67790 289128
rect 49602 288396 49608 288448
rect 49660 288436 49666 288448
rect 67634 288436 67640 288448
rect 49660 288408 67640 288436
rect 49660 288396 49666 288408
rect 67634 288396 67640 288408
rect 67692 288396 67698 288448
rect 67450 288328 67456 288380
rect 67508 288368 67514 288380
rect 67726 288368 67732 288380
rect 67508 288340 67732 288368
rect 67508 288328 67514 288340
rect 67726 288328 67732 288340
rect 67784 288328 67790 288380
rect 121454 288328 121460 288380
rect 121512 288368 121518 288380
rect 170398 288368 170404 288380
rect 121512 288340 170404 288368
rect 121512 288328 121518 288340
rect 170398 288328 170404 288340
rect 170456 288328 170462 288380
rect 172422 288328 172428 288380
rect 172480 288368 172486 288380
rect 176654 288368 176660 288380
rect 172480 288340 176660 288368
rect 172480 288328 172486 288340
rect 176654 288328 176660 288340
rect 176712 288328 176718 288380
rect 126422 287648 126428 287700
rect 126480 287688 126486 287700
rect 139394 287688 139400 287700
rect 126480 287660 139400 287688
rect 126480 287648 126486 287660
rect 139394 287648 139400 287660
rect 139452 287648 139458 287700
rect 50890 287036 50896 287088
rect 50948 287076 50954 287088
rect 67634 287076 67640 287088
rect 50948 287048 67640 287076
rect 50948 287036 50954 287048
rect 67634 287036 67640 287048
rect 67692 287036 67698 287088
rect 121638 287036 121644 287088
rect 121696 287076 121702 287088
rect 155218 287076 155224 287088
rect 121696 287048 155224 287076
rect 121696 287036 121702 287048
rect 155218 287036 155224 287048
rect 155276 287036 155282 287088
rect 131206 285744 131212 285796
rect 131264 285784 131270 285796
rect 132402 285784 132408 285796
rect 131264 285756 132408 285784
rect 131264 285744 131270 285756
rect 132402 285744 132408 285756
rect 132460 285784 132466 285796
rect 169386 285784 169392 285796
rect 132460 285756 169392 285784
rect 132460 285744 132466 285756
rect 169386 285744 169392 285756
rect 169444 285744 169450 285796
rect 54846 285676 54852 285728
rect 54904 285716 54910 285728
rect 67818 285716 67824 285728
rect 54904 285688 67824 285716
rect 54904 285676 54910 285688
rect 67818 285676 67824 285688
rect 67876 285676 67882 285728
rect 124398 285676 124404 285728
rect 124456 285716 124462 285728
rect 167914 285716 167920 285728
rect 124456 285688 167920 285716
rect 124456 285676 124462 285688
rect 167914 285676 167920 285688
rect 167972 285676 167978 285728
rect 295426 285676 295432 285728
rect 295484 285716 295490 285728
rect 308582 285716 308588 285728
rect 295484 285688 308588 285716
rect 295484 285676 295490 285688
rect 308582 285676 308588 285688
rect 308640 285676 308646 285728
rect 121546 285608 121552 285660
rect 121604 285648 121610 285660
rect 138014 285648 138020 285660
rect 121604 285620 138020 285648
rect 121604 285608 121610 285620
rect 138014 285608 138020 285620
rect 138072 285608 138078 285660
rect 121454 285540 121460 285592
rect 121512 285580 121518 285592
rect 131206 285580 131212 285592
rect 121512 285552 131212 285580
rect 121512 285540 121518 285552
rect 131206 285540 131212 285552
rect 131264 285540 131270 285592
rect 122190 284928 122196 284980
rect 122248 284968 122254 284980
rect 122834 284968 122840 284980
rect 122248 284940 122840 284968
rect 122248 284928 122254 284940
rect 122834 284928 122840 284940
rect 122892 284928 122898 284980
rect 130562 284928 130568 284980
rect 130620 284968 130626 284980
rect 156598 284968 156604 284980
rect 130620 284940 156604 284968
rect 130620 284928 130626 284940
rect 156598 284928 156604 284940
rect 156656 284928 156662 284980
rect 43990 284316 43996 284368
rect 44048 284356 44054 284368
rect 67634 284356 67640 284368
rect 44048 284328 67640 284356
rect 44048 284316 44054 284328
rect 67634 284316 67640 284328
rect 67692 284316 67698 284368
rect 53834 284248 53840 284300
rect 53892 284288 53898 284300
rect 67726 284288 67732 284300
rect 53892 284260 67732 284288
rect 53892 284248 53898 284260
rect 67726 284248 67732 284260
rect 67784 284248 67790 284300
rect 160830 284248 160836 284300
rect 160888 284288 160894 284300
rect 176654 284288 176660 284300
rect 160888 284260 176660 284288
rect 160888 284248 160894 284260
rect 176654 284248 176660 284260
rect 176712 284248 176718 284300
rect 66162 284180 66168 284232
rect 66220 284220 66226 284232
rect 67634 284220 67640 284232
rect 66220 284192 67640 284220
rect 66220 284180 66226 284192
rect 67634 284180 67640 284192
rect 67692 284180 67698 284232
rect 295426 283568 295432 283620
rect 295484 283608 295490 283620
rect 306558 283608 306564 283620
rect 295484 283580 306564 283608
rect 295484 283568 295490 283580
rect 306558 283568 306564 283580
rect 306616 283608 306622 283620
rect 325050 283608 325056 283620
rect 306616 283580 325056 283608
rect 306616 283568 306622 283580
rect 325050 283568 325056 283580
rect 325108 283568 325114 283620
rect 121454 282888 121460 282940
rect 121512 282928 121518 282940
rect 173250 282928 173256 282940
rect 121512 282900 173256 282928
rect 121512 282888 121518 282900
rect 173250 282888 173256 282900
rect 173308 282888 173314 282940
rect 123754 282820 123760 282872
rect 123812 282860 123818 282872
rect 166810 282860 166816 282872
rect 123812 282832 166816 282860
rect 123812 282820 123818 282832
rect 166810 282820 166816 282832
rect 166868 282860 166874 282872
rect 176654 282860 176660 282872
rect 166868 282832 176660 282860
rect 166868 282820 166874 282832
rect 176654 282820 176660 282832
rect 176712 282820 176718 282872
rect 121546 281596 121552 281648
rect 121604 281636 121610 281648
rect 152550 281636 152556 281648
rect 121604 281608 152556 281636
rect 121604 281596 121610 281608
rect 152550 281596 152556 281608
rect 152608 281596 152614 281648
rect 32950 281528 32956 281580
rect 33008 281568 33014 281580
rect 35710 281568 35716 281580
rect 33008 281540 35716 281568
rect 33008 281528 33014 281540
rect 35710 281528 35716 281540
rect 35768 281568 35774 281580
rect 35768 281540 67588 281568
rect 35768 281528 35774 281540
rect 67560 281500 67588 281540
rect 121454 281528 121460 281580
rect 121512 281568 121518 281580
rect 170398 281568 170404 281580
rect 121512 281540 170404 281568
rect 121512 281528 121518 281540
rect 170398 281528 170404 281540
rect 170456 281528 170462 281580
rect 295426 281528 295432 281580
rect 295484 281568 295490 281580
rect 359458 281568 359464 281580
rect 295484 281540 359464 281568
rect 295484 281528 295490 281540
rect 359458 281528 359464 281540
rect 359516 281528 359522 281580
rect 67634 281500 67640 281512
rect 67560 281472 67640 281500
rect 67634 281460 67640 281472
rect 67692 281460 67698 281512
rect 123662 280780 123668 280832
rect 123720 280820 123726 280832
rect 160094 280820 160100 280832
rect 123720 280792 160100 280820
rect 123720 280780 123726 280792
rect 160094 280780 160100 280792
rect 160152 280780 160158 280832
rect 55030 280168 55036 280220
rect 55088 280208 55094 280220
rect 67634 280208 67640 280220
rect 55088 280180 67640 280208
rect 55088 280168 55094 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121454 280168 121460 280220
rect 121512 280208 121518 280220
rect 136174 280208 136180 280220
rect 121512 280180 136180 280208
rect 121512 280168 121518 280180
rect 136174 280168 136180 280180
rect 136232 280168 136238 280220
rect 53742 280100 53748 280152
rect 53800 280140 53806 280152
rect 67726 280140 67732 280152
rect 53800 280112 67732 280140
rect 53800 280100 53806 280112
rect 67726 280100 67732 280112
rect 67784 280100 67790 280152
rect 169110 280100 169116 280152
rect 169168 280140 169174 280152
rect 176746 280140 176752 280152
rect 169168 280112 176752 280140
rect 169168 280100 169174 280112
rect 176746 280100 176752 280112
rect 176804 280100 176810 280152
rect 59078 280032 59084 280084
rect 59136 280072 59142 280084
rect 67634 280072 67640 280084
rect 59136 280044 67640 280072
rect 59136 280032 59142 280044
rect 67634 280032 67640 280044
rect 67692 280032 67698 280084
rect 22738 279420 22744 279472
rect 22796 279460 22802 279472
rect 59078 279460 59084 279472
rect 22796 279432 59084 279460
rect 22796 279420 22802 279432
rect 59078 279420 59084 279432
rect 59136 279420 59142 279472
rect 122742 279420 122748 279472
rect 122800 279460 122806 279472
rect 173158 279460 173164 279472
rect 122800 279432 173164 279460
rect 122800 279420 122806 279432
rect 173158 279420 173164 279432
rect 173216 279420 173222 279472
rect 295426 278808 295432 278860
rect 295484 278848 295490 278860
rect 297358 278848 297364 278860
rect 295484 278820 297364 278848
rect 295484 278808 295490 278820
rect 297358 278808 297364 278820
rect 297416 278808 297422 278860
rect 41230 278740 41236 278792
rect 41288 278780 41294 278792
rect 57238 278780 57244 278792
rect 41288 278752 57244 278780
rect 41288 278740 41294 278752
rect 57238 278740 57244 278752
rect 57296 278780 57302 278792
rect 57296 278752 57928 278780
rect 57296 278740 57302 278752
rect 57900 278712 57928 278752
rect 121454 278740 121460 278792
rect 121512 278780 121518 278792
rect 141418 278780 141424 278792
rect 121512 278752 141424 278780
rect 121512 278740 121518 278752
rect 141418 278740 141424 278752
rect 141476 278740 141482 278792
rect 67634 278712 67640 278724
rect 57900 278684 67640 278712
rect 67634 278672 67640 278684
rect 67692 278672 67698 278724
rect 121546 278672 121552 278724
rect 121604 278712 121610 278724
rect 129734 278712 129740 278724
rect 121604 278684 129740 278712
rect 121604 278672 121610 278684
rect 129734 278672 129740 278684
rect 129792 278672 129798 278724
rect 160094 278060 160100 278112
rect 160152 278100 160158 278112
rect 161382 278100 161388 278112
rect 160152 278072 161388 278100
rect 160152 278060 160158 278072
rect 161382 278060 161388 278072
rect 161440 278100 161446 278112
rect 176654 278100 176660 278112
rect 161440 278072 176660 278100
rect 161440 278060 161446 278072
rect 176654 278060 176660 278072
rect 176712 278060 176718 278112
rect 129734 277992 129740 278044
rect 129792 278032 129798 278044
rect 131022 278032 131028 278044
rect 129792 278004 131028 278032
rect 129792 277992 129798 278004
rect 131022 277992 131028 278004
rect 131080 278032 131086 278044
rect 169202 278032 169208 278044
rect 131080 278004 169208 278032
rect 131080 277992 131086 278004
rect 169202 277992 169208 278004
rect 169260 277992 169266 278044
rect 52178 277380 52184 277432
rect 52236 277420 52242 277432
rect 67634 277420 67640 277432
rect 52236 277392 67640 277420
rect 52236 277380 52242 277392
rect 67634 277380 67640 277392
rect 67692 277380 67698 277432
rect 145650 277420 145656 277432
rect 128280 277392 145656 277420
rect 121454 277312 121460 277364
rect 121512 277352 121518 277364
rect 127802 277352 127808 277364
rect 121512 277324 127808 277352
rect 121512 277312 121518 277324
rect 127802 277312 127808 277324
rect 127860 277352 127866 277364
rect 128280 277352 128308 277392
rect 145650 277380 145656 277392
rect 145708 277380 145714 277432
rect 127860 277324 128308 277352
rect 127860 277312 127866 277324
rect 62022 276088 62028 276140
rect 62080 276128 62086 276140
rect 64598 276128 64604 276140
rect 62080 276100 64604 276128
rect 62080 276088 62086 276100
rect 64598 276088 64604 276100
rect 64656 276128 64662 276140
rect 67634 276128 67640 276140
rect 64656 276100 67640 276128
rect 64656 276088 64662 276100
rect 67634 276088 67640 276100
rect 67692 276088 67698 276140
rect 50798 276020 50804 276072
rect 50856 276060 50862 276072
rect 67726 276060 67732 276072
rect 50856 276032 67732 276060
rect 50856 276020 50862 276032
rect 67726 276020 67732 276032
rect 67784 276020 67790 276072
rect 295426 276020 295432 276072
rect 295484 276060 295490 276072
rect 302418 276060 302424 276072
rect 295484 276032 302424 276060
rect 295484 276020 295490 276032
rect 302418 276020 302424 276032
rect 302476 276060 302482 276072
rect 306374 276060 306380 276072
rect 302476 276032 306380 276060
rect 302476 276020 302482 276032
rect 306374 276020 306380 276032
rect 306432 276020 306438 276072
rect 126514 275952 126520 276004
rect 126572 275992 126578 276004
rect 176654 275992 176660 276004
rect 126572 275964 176660 275992
rect 126572 275952 126578 275964
rect 176654 275952 176660 275964
rect 176712 275952 176718 276004
rect 65518 275476 65524 275528
rect 65576 275516 65582 275528
rect 68186 275516 68192 275528
rect 65576 275488 68192 275516
rect 65576 275476 65582 275488
rect 68186 275476 68192 275488
rect 68244 275476 68250 275528
rect 121454 274728 121460 274780
rect 121512 274768 121518 274780
rect 148594 274768 148600 274780
rect 121512 274740 148600 274768
rect 121512 274728 121518 274740
rect 148594 274728 148600 274740
rect 148652 274728 148658 274780
rect 49510 274660 49516 274712
rect 49568 274700 49574 274712
rect 67634 274700 67640 274712
rect 49568 274672 67640 274700
rect 49568 274660 49574 274672
rect 67634 274660 67640 274672
rect 67692 274660 67698 274712
rect 121546 274660 121552 274712
rect 121604 274700 121610 274712
rect 164970 274700 164976 274712
rect 121604 274672 164976 274700
rect 121604 274660 121610 274672
rect 164970 274660 164976 274672
rect 165028 274660 165034 274712
rect 295426 274660 295432 274712
rect 295484 274700 295490 274712
rect 301130 274700 301136 274712
rect 295484 274672 301136 274700
rect 295484 274660 295490 274672
rect 301130 274660 301136 274672
rect 301188 274660 301194 274712
rect 39942 274592 39948 274644
rect 40000 274632 40006 274644
rect 68002 274632 68008 274644
rect 40000 274604 68008 274632
rect 40000 274592 40006 274604
rect 68002 274592 68008 274604
rect 68060 274592 68066 274644
rect 121454 274592 121460 274644
rect 121512 274632 121518 274644
rect 179874 274632 179880 274644
rect 121512 274604 179880 274632
rect 121512 274592 121518 274604
rect 179874 274592 179880 274604
rect 179932 274592 179938 274644
rect 65978 273232 65984 273284
rect 66036 273272 66042 273284
rect 67818 273272 67824 273284
rect 66036 273244 67824 273272
rect 66036 273232 66042 273244
rect 67818 273232 67824 273244
rect 67876 273232 67882 273284
rect 121454 273232 121460 273284
rect 121512 273272 121518 273284
rect 158070 273272 158076 273284
rect 121512 273244 158076 273272
rect 121512 273232 121518 273244
rect 158070 273232 158076 273244
rect 158128 273232 158134 273284
rect 295426 272688 295432 272740
rect 295484 272728 295490 272740
rect 298278 272728 298284 272740
rect 295484 272700 298284 272728
rect 295484 272688 295490 272700
rect 298278 272688 298284 272700
rect 298336 272688 298342 272740
rect 121454 272552 121460 272604
rect 121512 272592 121518 272604
rect 124214 272592 124220 272604
rect 121512 272564 124220 272592
rect 121512 272552 121518 272564
rect 124214 272552 124220 272564
rect 124272 272592 124278 272604
rect 147122 272592 147128 272604
rect 124272 272564 147128 272592
rect 124272 272552 124278 272564
rect 147122 272552 147128 272564
rect 147180 272552 147186 272604
rect 128354 272484 128360 272536
rect 128412 272524 128418 272536
rect 129274 272524 129280 272536
rect 128412 272496 129280 272524
rect 128412 272484 128418 272496
rect 129274 272484 129280 272496
rect 129332 272524 129338 272536
rect 176654 272524 176660 272536
rect 129332 272496 176660 272524
rect 129332 272484 129338 272496
rect 176654 272484 176660 272496
rect 176712 272484 176718 272536
rect 66162 271940 66168 271992
rect 66220 271980 66226 271992
rect 67818 271980 67824 271992
rect 66220 271952 67824 271980
rect 66220 271940 66226 271952
rect 67818 271940 67824 271952
rect 67876 271940 67882 271992
rect 57790 271872 57796 271924
rect 57848 271912 57854 271924
rect 67634 271912 67640 271924
rect 57848 271884 67640 271912
rect 57848 271872 57854 271884
rect 67634 271872 67640 271884
rect 67692 271872 67698 271924
rect 61838 270580 61844 270632
rect 61896 270620 61902 270632
rect 67634 270620 67640 270632
rect 61896 270592 67640 270620
rect 61896 270580 61902 270592
rect 67634 270580 67640 270592
rect 67692 270580 67698 270632
rect 56318 270512 56324 270564
rect 56376 270552 56382 270564
rect 67726 270552 67732 270564
rect 56376 270524 67732 270552
rect 56376 270512 56382 270524
rect 67726 270512 67732 270524
rect 67784 270512 67790 270564
rect 121454 270512 121460 270564
rect 121512 270552 121518 270564
rect 138750 270552 138756 270564
rect 121512 270524 138756 270552
rect 121512 270512 121518 270524
rect 138750 270512 138756 270524
rect 138808 270512 138814 270564
rect 54938 269764 54944 269816
rect 54996 269804 55002 269816
rect 67634 269804 67640 269816
rect 54996 269776 67640 269804
rect 54996 269764 55002 269776
rect 67634 269764 67640 269776
rect 67692 269764 67698 269816
rect 120902 269764 120908 269816
rect 120960 269804 120966 269816
rect 128354 269804 128360 269816
rect 120960 269776 128360 269804
rect 120960 269764 120966 269776
rect 128354 269764 128360 269776
rect 128412 269764 128418 269816
rect 121454 269152 121460 269204
rect 121512 269192 121518 269204
rect 154022 269192 154028 269204
rect 121512 269164 154028 269192
rect 121512 269152 121518 269164
rect 154022 269152 154028 269164
rect 154080 269152 154086 269204
rect 62022 269084 62028 269136
rect 62080 269124 62086 269136
rect 67726 269124 67732 269136
rect 62080 269096 67732 269124
rect 62080 269084 62086 269096
rect 67726 269084 67732 269096
rect 67784 269084 67790 269136
rect 121546 269084 121552 269136
rect 121604 269124 121610 269136
rect 160830 269124 160836 269136
rect 121604 269096 160836 269124
rect 121604 269084 121610 269096
rect 160830 269084 160836 269096
rect 160888 269084 160894 269136
rect 295426 269084 295432 269136
rect 295484 269124 295490 269136
rect 349338 269124 349344 269136
rect 295484 269096 349344 269124
rect 295484 269084 295490 269096
rect 349338 269084 349344 269096
rect 349396 269084 349402 269136
rect 121454 269016 121460 269068
rect 121512 269056 121518 269068
rect 135990 269056 135996 269068
rect 121512 269028 135996 269056
rect 121512 269016 121518 269028
rect 135990 269016 135996 269028
rect 136048 269016 136054 269068
rect 121454 268336 121460 268388
rect 121512 268376 121518 268388
rect 126238 268376 126244 268388
rect 121512 268348 126244 268376
rect 121512 268336 121518 268348
rect 126238 268336 126244 268348
rect 126296 268336 126302 268388
rect 64782 267792 64788 267844
rect 64840 267832 64846 267844
rect 67726 267832 67732 267844
rect 64840 267804 67732 267832
rect 64840 267792 64846 267804
rect 67726 267792 67732 267804
rect 67784 267792 67790 267844
rect 46750 267724 46756 267776
rect 46808 267764 46814 267776
rect 67634 267764 67640 267776
rect 46808 267736 67640 267764
rect 46808 267724 46814 267736
rect 67634 267724 67640 267736
rect 67692 267724 67698 267776
rect 121546 267656 121552 267708
rect 121604 267696 121610 267708
rect 148318 267696 148324 267708
rect 121604 267668 148324 267696
rect 121604 267656 121610 267668
rect 148318 267656 148324 267668
rect 148376 267656 148382 267708
rect 3418 266976 3424 267028
rect 3476 267016 3482 267028
rect 13078 267016 13084 267028
rect 3476 266988 13084 267016
rect 3476 266976 3482 266988
rect 13078 266976 13084 266988
rect 13136 266976 13142 267028
rect 121454 266364 121460 266416
rect 121512 266404 121518 266416
rect 166350 266404 166356 266416
rect 121512 266376 166356 266404
rect 121512 266364 121518 266376
rect 166350 266364 166356 266376
rect 166408 266364 166414 266416
rect 49418 266296 49424 266348
rect 49476 266336 49482 266348
rect 67634 266336 67640 266348
rect 49476 266308 67640 266336
rect 49476 266296 49482 266308
rect 67634 266296 67640 266308
rect 67692 266296 67698 266348
rect 53466 264936 53472 264988
rect 53524 264976 53530 264988
rect 68094 264976 68100 264988
rect 53524 264948 68100 264976
rect 53524 264936 53530 264948
rect 68094 264936 68100 264948
rect 68152 264936 68158 264988
rect 295426 264936 295432 264988
rect 295484 264976 295490 264988
rect 325050 264976 325056 264988
rect 295484 264948 325056 264976
rect 295484 264936 295490 264948
rect 325050 264936 325056 264948
rect 325108 264936 325114 264988
rect 121454 264188 121460 264240
rect 121512 264228 121518 264240
rect 159358 264228 159364 264240
rect 121512 264200 159364 264228
rect 121512 264188 121518 264200
rect 159358 264188 159364 264200
rect 159416 264188 159422 264240
rect 18598 263576 18604 263628
rect 18656 263616 18662 263628
rect 59078 263616 59084 263628
rect 18656 263588 59084 263616
rect 18656 263576 18662 263588
rect 59078 263576 59084 263588
rect 59136 263616 59142 263628
rect 67634 263616 67640 263628
rect 59136 263588 67640 263616
rect 59136 263576 59142 263588
rect 67634 263576 67640 263588
rect 67692 263576 67698 263628
rect 121546 263576 121552 263628
rect 121604 263616 121610 263628
rect 146938 263616 146944 263628
rect 121604 263588 146944 263616
rect 121604 263576 121610 263588
rect 146938 263576 146944 263588
rect 146996 263576 147002 263628
rect 121454 263508 121460 263560
rect 121512 263548 121518 263560
rect 129826 263548 129832 263560
rect 121512 263520 129832 263548
rect 121512 263508 121518 263520
rect 129826 263508 129832 263520
rect 129884 263508 129890 263560
rect 4062 262828 4068 262880
rect 4120 262868 4126 262880
rect 62114 262868 62120 262880
rect 4120 262840 62120 262868
rect 4120 262828 4126 262840
rect 62114 262828 62120 262840
rect 62172 262828 62178 262880
rect 121454 262828 121460 262880
rect 121512 262868 121518 262880
rect 124306 262868 124312 262880
rect 121512 262840 124312 262868
rect 121512 262828 121518 262840
rect 124306 262828 124312 262840
rect 124364 262868 124370 262880
rect 140222 262868 140228 262880
rect 124364 262840 140228 262868
rect 124364 262828 124370 262840
rect 140222 262828 140228 262840
rect 140280 262828 140286 262880
rect 63310 262284 63316 262336
rect 63368 262324 63374 262336
rect 67726 262324 67732 262336
rect 63368 262296 67732 262324
rect 63368 262284 63374 262296
rect 67726 262284 67732 262296
rect 67784 262284 67790 262336
rect 53742 262216 53748 262268
rect 53800 262256 53806 262268
rect 67634 262256 67640 262268
rect 53800 262228 67640 262256
rect 53800 262216 53806 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 120718 262216 120724 262268
rect 120776 262256 120782 262268
rect 120994 262256 121000 262268
rect 120776 262228 121000 262256
rect 120776 262216 120782 262228
rect 120994 262216 121000 262228
rect 121052 262256 121058 262268
rect 167730 262256 167736 262268
rect 121052 262228 167736 262256
rect 121052 262216 121058 262228
rect 167730 262216 167736 262228
rect 167788 262216 167794 262268
rect 62206 262148 62212 262200
rect 62264 262188 62270 262200
rect 63034 262188 63040 262200
rect 62264 262160 63040 262188
rect 62264 262148 62270 262160
rect 63034 262148 63040 262160
rect 63092 262188 63098 262200
rect 67726 262188 67732 262200
rect 63092 262160 67732 262188
rect 63092 262148 63098 262160
rect 67726 262148 67732 262160
rect 67784 262148 67790 262200
rect 121454 262148 121460 262200
rect 121512 262188 121518 262200
rect 171962 262188 171968 262200
rect 121512 262160 171968 262188
rect 121512 262148 121518 262160
rect 171962 262148 171968 262160
rect 172020 262148 172026 262200
rect 140130 262080 140136 262132
rect 140188 262120 140194 262132
rect 176654 262120 176660 262132
rect 140188 262092 176660 262120
rect 140188 262080 140194 262092
rect 176654 262080 176660 262092
rect 176712 262080 176718 262132
rect 61746 261536 61752 261588
rect 61804 261576 61810 261588
rect 61930 261576 61936 261588
rect 61804 261548 61936 261576
rect 61804 261536 61810 261548
rect 61930 261536 61936 261548
rect 61988 261576 61994 261588
rect 67634 261576 67640 261588
rect 61988 261548 67640 261576
rect 61988 261536 61994 261548
rect 67634 261536 67640 261548
rect 67692 261536 67698 261588
rect 50706 261468 50712 261520
rect 50764 261508 50770 261520
rect 62206 261508 62212 261520
rect 50764 261480 62212 261508
rect 50764 261468 50770 261480
rect 62206 261468 62212 261480
rect 62264 261468 62270 261520
rect 52270 260856 52276 260908
rect 52328 260896 52334 260908
rect 52328 260868 55214 260896
rect 52328 260856 52334 260868
rect 55186 260828 55214 260868
rect 295426 260856 295432 260908
rect 295484 260896 295490 260908
rect 309686 260896 309692 260908
rect 295484 260868 309692 260896
rect 295484 260856 295490 260868
rect 309686 260856 309692 260868
rect 309744 260856 309750 260908
rect 55858 260828 55864 260840
rect 55186 260800 55864 260828
rect 55858 260788 55864 260800
rect 55916 260828 55922 260840
rect 67726 260828 67732 260840
rect 55916 260800 67732 260828
rect 55916 260788 55922 260800
rect 67726 260788 67732 260800
rect 67784 260788 67790 260840
rect 121454 260788 121460 260840
rect 121512 260828 121518 260840
rect 161474 260828 161480 260840
rect 121512 260800 161480 260828
rect 121512 260788 121518 260800
rect 161474 260788 161480 260800
rect 161532 260788 161538 260840
rect 62114 260720 62120 260772
rect 62172 260760 62178 260772
rect 67634 260760 67640 260772
rect 62172 260732 67640 260760
rect 62172 260720 62178 260732
rect 67634 260720 67640 260732
rect 67692 260720 67698 260772
rect 122098 260108 122104 260160
rect 122156 260148 122162 260160
rect 141602 260148 141608 260160
rect 122156 260120 141608 260148
rect 122156 260108 122162 260120
rect 141602 260108 141608 260120
rect 141660 260108 141666 260160
rect 121454 259428 121460 259480
rect 121512 259468 121518 259480
rect 160922 259468 160928 259480
rect 121512 259440 160928 259468
rect 121512 259428 121518 259440
rect 160922 259428 160928 259440
rect 160980 259428 160986 259480
rect 347038 259360 347044 259412
rect 347096 259400 347102 259412
rect 580166 259400 580172 259412
rect 347096 259372 580172 259400
rect 347096 259360 347102 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 122282 258680 122288 258732
rect 122340 258720 122346 258732
rect 171962 258720 171968 258732
rect 122340 258692 171968 258720
rect 122340 258680 122346 258692
rect 171962 258680 171968 258692
rect 172020 258680 172026 258732
rect 57698 258136 57704 258188
rect 57756 258176 57762 258188
rect 67634 258176 67640 258188
rect 57756 258148 67640 258176
rect 57756 258136 57762 258148
rect 67634 258136 67640 258148
rect 67692 258136 67698 258188
rect 56410 258068 56416 258120
rect 56468 258108 56474 258120
rect 67726 258108 67732 258120
rect 56468 258080 67732 258108
rect 56468 258068 56474 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 121454 258068 121460 258120
rect 121512 258108 121518 258120
rect 162302 258108 162308 258120
rect 121512 258080 162308 258108
rect 121512 258068 121518 258080
rect 162302 258068 162308 258080
rect 162360 258068 162366 258120
rect 52086 258000 52092 258052
rect 52144 258040 52150 258052
rect 67634 258040 67640 258052
rect 52144 258012 67640 258040
rect 52144 258000 52150 258012
rect 67634 258000 67640 258012
rect 67692 258000 67698 258052
rect 14458 257320 14464 257372
rect 14516 257360 14522 257372
rect 52086 257360 52092 257372
rect 14516 257332 52092 257360
rect 14516 257320 14522 257332
rect 52086 257320 52092 257332
rect 52144 257320 52150 257372
rect 170950 257320 170956 257372
rect 171008 257360 171014 257372
rect 178678 257360 178684 257372
rect 171008 257332 178684 257360
rect 171008 257320 171014 257332
rect 178678 257320 178684 257332
rect 178736 257320 178742 257372
rect 121546 256844 121552 256896
rect 121604 256884 121610 256896
rect 148318 256884 148324 256896
rect 121604 256856 148324 256884
rect 121604 256844 121610 256856
rect 148318 256844 148324 256856
rect 148376 256844 148382 256896
rect 121454 256776 121460 256828
rect 121512 256816 121518 256828
rect 156598 256816 156604 256828
rect 121512 256788 156604 256816
rect 121512 256776 121518 256788
rect 156598 256776 156604 256788
rect 156656 256776 156662 256828
rect 123570 256708 123576 256760
rect 123628 256748 123634 256760
rect 176654 256748 176660 256760
rect 123628 256720 176660 256748
rect 123628 256708 123634 256720
rect 176654 256708 176660 256720
rect 176712 256708 176718 256760
rect 59262 255960 59268 256012
rect 59320 256000 59326 256012
rect 67910 256000 67916 256012
rect 59320 255972 67916 256000
rect 59320 255960 59326 255972
rect 67910 255960 67916 255972
rect 67968 255960 67974 256012
rect 122466 255960 122472 256012
rect 122524 256000 122530 256012
rect 130378 256000 130384 256012
rect 122524 255972 130384 256000
rect 122524 255960 122530 255972
rect 130378 255960 130384 255972
rect 130436 255960 130442 256012
rect 121546 255348 121552 255400
rect 121604 255388 121610 255400
rect 135162 255388 135168 255400
rect 121604 255360 135168 255388
rect 121604 255348 121610 255360
rect 135162 255348 135168 255360
rect 135220 255388 135226 255400
rect 140774 255388 140780 255400
rect 135220 255360 140780 255388
rect 135220 255348 135226 255360
rect 140774 255348 140780 255360
rect 140832 255348 140838 255400
rect 60550 255280 60556 255332
rect 60608 255320 60614 255332
rect 67634 255320 67640 255332
rect 60608 255292 67640 255320
rect 60608 255280 60614 255292
rect 67634 255280 67640 255292
rect 67692 255280 67698 255332
rect 121454 255280 121460 255332
rect 121512 255320 121518 255332
rect 162394 255320 162400 255332
rect 121512 255292 162400 255320
rect 121512 255280 121518 255292
rect 162394 255280 162400 255292
rect 162452 255280 162458 255332
rect 41322 255212 41328 255264
rect 41380 255252 41386 255264
rect 62114 255252 62120 255264
rect 41380 255224 62120 255252
rect 41380 255212 41386 255224
rect 62114 255212 62120 255224
rect 62172 255212 62178 255264
rect 62114 254532 62120 254584
rect 62172 254572 62178 254584
rect 63126 254572 63132 254584
rect 62172 254544 63132 254572
rect 62172 254532 62178 254544
rect 63126 254532 63132 254544
rect 63184 254572 63190 254584
rect 67634 254572 67640 254584
rect 63184 254544 67640 254572
rect 63184 254532 63190 254544
rect 67634 254532 67640 254544
rect 67692 254532 67698 254584
rect 121454 253988 121460 254040
rect 121512 254028 121518 254040
rect 151262 254028 151268 254040
rect 121512 254000 151268 254028
rect 121512 253988 121518 254000
rect 151262 253988 151268 254000
rect 151320 253988 151326 254040
rect 3418 253920 3424 253972
rect 3476 253960 3482 253972
rect 26878 253960 26884 253972
rect 3476 253932 26884 253960
rect 3476 253920 3482 253932
rect 26878 253920 26884 253932
rect 26936 253920 26942 253972
rect 61930 253920 61936 253972
rect 61988 253960 61994 253972
rect 67726 253960 67732 253972
rect 61988 253932 67732 253960
rect 61988 253920 61994 253932
rect 67726 253920 67732 253932
rect 67784 253920 67790 253972
rect 120718 253920 120724 253972
rect 120776 253960 120782 253972
rect 172330 253960 172336 253972
rect 120776 253932 172336 253960
rect 120776 253920 120782 253932
rect 172330 253920 172336 253932
rect 172388 253960 172394 253972
rect 176654 253960 176660 253972
rect 172388 253932 176660 253960
rect 172388 253920 172394 253932
rect 176654 253920 176660 253932
rect 176712 253920 176718 253972
rect 295518 253920 295524 253972
rect 295576 253960 295582 253972
rect 311158 253960 311164 253972
rect 295576 253932 311164 253960
rect 295576 253920 295582 253932
rect 311158 253920 311164 253932
rect 311216 253920 311222 253972
rect 62114 253852 62120 253904
rect 62172 253892 62178 253904
rect 62758 253892 62764 253904
rect 62172 253864 62764 253892
rect 62172 253852 62178 253864
rect 62758 253852 62764 253864
rect 62816 253892 62822 253904
rect 67634 253892 67640 253904
rect 62816 253864 67640 253892
rect 62816 253852 62822 253864
rect 67634 253852 67640 253864
rect 67692 253852 67698 253904
rect 121454 253852 121460 253904
rect 121512 253892 121518 253904
rect 166258 253892 166264 253904
rect 121512 253864 166264 253892
rect 121512 253852 121518 253864
rect 166258 253852 166264 253864
rect 166316 253852 166322 253904
rect 21358 253172 21364 253224
rect 21416 253212 21422 253224
rect 62114 253212 62120 253224
rect 21416 253184 62120 253212
rect 21416 253172 21422 253184
rect 62114 253172 62120 253184
rect 62172 253172 62178 253224
rect 121546 252560 121552 252612
rect 121604 252600 121610 252612
rect 138842 252600 138848 252612
rect 121604 252572 138848 252600
rect 121604 252560 121610 252572
rect 138842 252560 138848 252572
rect 138900 252560 138906 252612
rect 166718 252560 166724 252612
rect 166776 252600 166782 252612
rect 176654 252600 176660 252612
rect 166776 252572 176660 252600
rect 166776 252560 166782 252572
rect 176654 252560 176660 252572
rect 176712 252560 176718 252612
rect 62114 251812 62120 251864
rect 62172 251852 62178 251864
rect 63402 251852 63408 251864
rect 62172 251824 63408 251852
rect 62172 251812 62178 251824
rect 63402 251812 63408 251824
rect 63460 251852 63466 251864
rect 67634 251852 67640 251864
rect 63460 251824 67640 251852
rect 63460 251812 63466 251824
rect 67634 251812 67640 251824
rect 67692 251812 67698 251864
rect 295518 251812 295524 251864
rect 295576 251852 295582 251864
rect 298370 251852 298376 251864
rect 295576 251824 298376 251852
rect 295576 251812 295582 251824
rect 298370 251812 298376 251824
rect 298428 251852 298434 251864
rect 304994 251852 305000 251864
rect 298428 251824 305000 251852
rect 298428 251812 298434 251824
rect 304994 251812 305000 251824
rect 305052 251812 305058 251864
rect 45186 251200 45192 251252
rect 45244 251240 45250 251252
rect 62114 251240 62120 251252
rect 45244 251212 62120 251240
rect 45244 251200 45250 251212
rect 62114 251200 62120 251212
rect 62172 251200 62178 251252
rect 121454 251200 121460 251252
rect 121512 251240 121518 251252
rect 176102 251240 176108 251252
rect 121512 251212 176108 251240
rect 121512 251200 121518 251212
rect 176102 251200 176108 251212
rect 176160 251200 176166 251252
rect 120626 251132 120632 251184
rect 120684 251172 120690 251184
rect 133966 251172 133972 251184
rect 120684 251144 133972 251172
rect 120684 251132 120690 251144
rect 133966 251132 133972 251144
rect 134024 251132 134030 251184
rect 58710 249840 58716 249892
rect 58768 249880 58774 249892
rect 67634 249880 67640 249892
rect 58768 249852 67640 249880
rect 58768 249840 58774 249852
rect 67634 249840 67640 249852
rect 67692 249840 67698 249892
rect 121546 249772 121552 249824
rect 121604 249812 121610 249824
rect 134518 249812 134524 249824
rect 121604 249784 134524 249812
rect 121604 249772 121610 249784
rect 134518 249772 134524 249784
rect 134576 249772 134582 249824
rect 166810 249772 166816 249824
rect 166868 249812 166874 249824
rect 176654 249812 176660 249824
rect 166868 249784 176660 249812
rect 166868 249772 166874 249784
rect 176654 249772 176660 249784
rect 176712 249772 176718 249824
rect 295518 249772 295524 249824
rect 295576 249812 295582 249824
rect 325142 249812 325148 249824
rect 295576 249784 325148 249812
rect 295576 249772 295582 249784
rect 325142 249772 325148 249784
rect 325200 249772 325206 249824
rect 45462 249704 45468 249756
rect 45520 249744 45526 249756
rect 67634 249744 67640 249756
rect 45520 249716 67640 249744
rect 45520 249704 45526 249716
rect 67634 249704 67640 249716
rect 67692 249704 67698 249756
rect 121454 249704 121460 249756
rect 121512 249744 121518 249756
rect 130470 249744 130476 249756
rect 121512 249716 130476 249744
rect 121512 249704 121518 249716
rect 130470 249704 130476 249716
rect 130528 249704 130534 249756
rect 48222 249636 48228 249688
rect 48280 249676 48286 249688
rect 58710 249676 58716 249688
rect 48280 249648 58716 249676
rect 48280 249636 48286 249648
rect 58710 249636 58716 249648
rect 58768 249636 58774 249688
rect 63126 248412 63132 248464
rect 63184 248452 63190 248464
rect 67634 248452 67640 248464
rect 63184 248424 67640 248452
rect 63184 248412 63190 248424
rect 67634 248412 67640 248424
rect 67692 248412 67698 248464
rect 121454 248344 121460 248396
rect 121512 248384 121518 248396
rect 174538 248384 174544 248396
rect 121512 248356 174544 248384
rect 121512 248344 121518 248356
rect 174538 248344 174544 248356
rect 174596 248344 174602 248396
rect 64690 247120 64696 247172
rect 64748 247160 64754 247172
rect 67634 247160 67640 247172
rect 64748 247132 67640 247160
rect 64748 247120 64754 247132
rect 67634 247120 67640 247132
rect 67692 247120 67698 247172
rect 63218 247052 63224 247104
rect 63276 247092 63282 247104
rect 67726 247092 67732 247104
rect 63276 247064 67732 247092
rect 63276 247052 63282 247064
rect 67726 247052 67732 247064
rect 67784 247052 67790 247104
rect 121546 247052 121552 247104
rect 121604 247092 121610 247104
rect 144362 247092 144368 247104
rect 121604 247064 144368 247092
rect 121604 247052 121610 247064
rect 144362 247052 144368 247064
rect 144420 247052 144426 247104
rect 50982 246984 50988 247036
rect 51040 247024 51046 247036
rect 67634 247024 67640 247036
rect 51040 246996 67640 247024
rect 51040 246984 51046 246996
rect 67634 246984 67640 246996
rect 67692 246984 67698 247036
rect 128354 246984 128360 247036
rect 128412 247024 128418 247036
rect 132494 247024 132500 247036
rect 128412 246996 132500 247024
rect 128412 246984 128418 246996
rect 132494 246984 132500 246996
rect 132552 247024 132558 247036
rect 176654 247024 176660 247036
rect 132552 246996 176660 247024
rect 132552 246984 132558 246996
rect 176654 246984 176660 246996
rect 176712 246984 176718 247036
rect 66070 246916 66076 246968
rect 66128 246956 66134 246968
rect 68186 246956 68192 246968
rect 66128 246928 68192 246956
rect 66128 246916 66134 246928
rect 68186 246916 68192 246928
rect 68244 246916 68250 246968
rect 139302 245760 139308 245812
rect 139360 245800 139366 245812
rect 140130 245800 140136 245812
rect 139360 245772 140136 245800
rect 139360 245760 139366 245772
rect 140130 245760 140136 245772
rect 140188 245760 140194 245812
rect 121546 245692 121552 245744
rect 121604 245732 121610 245744
rect 147030 245732 147036 245744
rect 121604 245704 147036 245732
rect 121604 245692 121610 245704
rect 147030 245692 147036 245704
rect 147088 245692 147094 245744
rect 121454 245624 121460 245676
rect 121512 245664 121518 245676
rect 152642 245664 152648 245676
rect 121512 245636 152648 245664
rect 121512 245624 121518 245636
rect 152642 245624 152648 245636
rect 152700 245624 152706 245676
rect 295518 245624 295524 245676
rect 295576 245664 295582 245676
rect 512638 245664 512644 245676
rect 295576 245636 512644 245664
rect 295576 245624 295582 245636
rect 512638 245624 512644 245636
rect 512696 245624 512702 245676
rect 121546 245556 121552 245608
rect 121604 245596 121610 245608
rect 164234 245596 164240 245608
rect 121604 245568 164240 245596
rect 121604 245556 121610 245568
rect 164234 245556 164240 245568
rect 164292 245556 164298 245608
rect 121454 245012 121460 245064
rect 121512 245052 121518 245064
rect 140130 245052 140136 245064
rect 121512 245024 140136 245052
rect 121512 245012 121518 245024
rect 140130 245012 140136 245024
rect 140188 245012 140194 245064
rect 134610 244944 134616 244996
rect 134668 244984 134674 244996
rect 164878 244984 164884 244996
rect 134668 244956 164884 244984
rect 134668 244944 134674 244956
rect 164878 244944 164884 244956
rect 164936 244944 164942 244996
rect 120810 244876 120816 244928
rect 120868 244916 120874 244928
rect 172054 244916 172060 244928
rect 120868 244888 172060 244916
rect 120868 244876 120874 244888
rect 172054 244876 172060 244888
rect 172112 244876 172118 244928
rect 66070 244264 66076 244316
rect 66128 244304 66134 244316
rect 68186 244304 68192 244316
rect 66128 244276 68192 244304
rect 66128 244264 66134 244276
rect 68186 244264 68192 244276
rect 68244 244264 68250 244316
rect 8938 244196 8944 244248
rect 8996 244236 9002 244248
rect 39666 244236 39672 244248
rect 8996 244208 39672 244236
rect 8996 244196 9002 244208
rect 39666 244196 39672 244208
rect 39724 244236 39730 244248
rect 67634 244236 67640 244248
rect 39724 244208 67640 244236
rect 39724 244196 39730 244208
rect 67634 244196 67640 244208
rect 67692 244196 67698 244248
rect 121454 244196 121460 244248
rect 121512 244236 121518 244248
rect 153838 244236 153844 244248
rect 121512 244208 153844 244236
rect 121512 244196 121518 244208
rect 153838 244196 153844 244208
rect 153896 244196 153902 244248
rect 296898 242904 296904 242956
rect 296956 242944 296962 242956
rect 347038 242944 347044 242956
rect 296956 242916 347044 242944
rect 296956 242904 296962 242916
rect 347038 242904 347044 242916
rect 347096 242904 347102 242956
rect 34422 242836 34428 242888
rect 34480 242876 34486 242888
rect 69658 242876 69664 242888
rect 34480 242848 69664 242876
rect 34480 242836 34486 242848
rect 69658 242836 69664 242848
rect 69716 242836 69722 242888
rect 121546 242836 121552 242888
rect 121604 242876 121610 242888
rect 143534 242876 143540 242888
rect 121604 242848 143540 242876
rect 121604 242836 121610 242848
rect 143534 242836 143540 242848
rect 143592 242836 143598 242888
rect 64598 242768 64604 242820
rect 64656 242808 64662 242820
rect 66990 242808 66996 242820
rect 64656 242780 66996 242808
rect 64656 242768 64662 242780
rect 66990 242768 66996 242780
rect 67048 242768 67054 242820
rect 121454 242768 121460 242820
rect 121512 242808 121518 242820
rect 127710 242808 127716 242820
rect 121512 242780 127716 242808
rect 121512 242768 121518 242780
rect 127710 242768 127716 242780
rect 127768 242768 127774 242820
rect 119982 242224 119988 242276
rect 120040 242264 120046 242276
rect 155954 242264 155960 242276
rect 120040 242236 155960 242264
rect 120040 242224 120046 242236
rect 155954 242224 155960 242236
rect 156012 242224 156018 242276
rect 119890 242156 119896 242208
rect 119948 242196 119954 242208
rect 179414 242196 179420 242208
rect 119948 242168 179420 242196
rect 119948 242156 119954 242168
rect 179414 242156 179420 242168
rect 179472 242156 179478 242208
rect 63402 241544 63408 241596
rect 63460 241584 63466 241596
rect 67634 241584 67640 241596
rect 63460 241556 67640 241584
rect 63460 241544 63466 241556
rect 67634 241544 67640 241556
rect 67692 241544 67698 241596
rect 60458 241476 60464 241528
rect 60516 241516 60522 241528
rect 67726 241516 67732 241528
rect 60516 241488 67732 241516
rect 60516 241476 60522 241488
rect 67726 241476 67732 241488
rect 67784 241476 67790 241528
rect 53558 241408 53564 241460
rect 53616 241448 53622 241460
rect 67634 241448 67640 241460
rect 53616 241420 67640 241448
rect 53616 241408 53622 241420
rect 67634 241408 67640 241420
rect 67692 241408 67698 241460
rect 155310 241408 155316 241460
rect 155368 241448 155374 241460
rect 298278 241448 298284 241460
rect 155368 241420 298284 241448
rect 155368 241408 155374 241420
rect 298278 241408 298284 241420
rect 298336 241408 298342 241460
rect 42702 240728 42708 240780
rect 42760 240768 42766 240780
rect 63586 240768 63592 240780
rect 42760 240740 63592 240768
rect 42760 240728 42766 240740
rect 63586 240728 63592 240740
rect 63644 240728 63650 240780
rect 135162 240728 135168 240780
rect 135220 240768 135226 240780
rect 135220 240740 180794 240768
rect 135220 240728 135226 240740
rect 180766 240632 180794 240740
rect 189994 240632 190000 240644
rect 180766 240604 190000 240632
rect 189994 240592 190000 240604
rect 190052 240592 190058 240644
rect 292022 240592 292028 240644
rect 292080 240632 292086 240644
rect 293310 240632 293316 240644
rect 292080 240604 293316 240632
rect 292080 240592 292086 240604
rect 293310 240592 293316 240604
rect 293368 240592 293374 240644
rect 63586 240116 63592 240168
rect 63644 240156 63650 240168
rect 64598 240156 64604 240168
rect 63644 240128 64604 240156
rect 63644 240116 63650 240128
rect 64598 240116 64604 240128
rect 64656 240156 64662 240168
rect 67634 240156 67640 240168
rect 64656 240128 67640 240156
rect 64656 240116 64662 240128
rect 67634 240116 67640 240128
rect 67692 240116 67698 240168
rect 121454 240116 121460 240168
rect 121512 240156 121518 240168
rect 153838 240156 153844 240168
rect 121512 240128 153844 240156
rect 121512 240116 121518 240128
rect 153838 240116 153844 240128
rect 153896 240116 153902 240168
rect 163590 240048 163596 240100
rect 163648 240088 163654 240100
rect 580166 240088 580172 240100
rect 163648 240060 580172 240088
rect 163648 240048 163654 240060
rect 580166 240048 580172 240060
rect 580224 240048 580230 240100
rect 121546 239980 121552 240032
rect 121604 240020 121610 240032
rect 309134 240020 309140 240032
rect 121604 239992 309140 240020
rect 121604 239980 121610 239992
rect 309134 239980 309140 239992
rect 309192 240020 309198 240032
rect 310422 240020 310428 240032
rect 309192 239992 310428 240020
rect 309192 239980 309198 239992
rect 310422 239980 310428 239992
rect 310480 239980 310486 240032
rect 66254 239912 66260 239964
rect 66312 239952 66318 239964
rect 70670 239952 70676 239964
rect 66312 239924 70676 239952
rect 66312 239912 66318 239924
rect 70670 239912 70676 239924
rect 70728 239912 70734 239964
rect 118970 239912 118976 239964
rect 119028 239952 119034 239964
rect 119890 239952 119896 239964
rect 119028 239924 119896 239952
rect 119028 239912 119034 239924
rect 119890 239912 119896 239924
rect 119948 239912 119954 239964
rect 156598 239912 156604 239964
rect 156656 239952 156662 239964
rect 306558 239952 306564 239964
rect 156656 239924 306564 239952
rect 156656 239912 156662 239924
rect 306558 239912 306564 239924
rect 306616 239912 306622 239964
rect 117038 239844 117044 239896
rect 117096 239884 117102 239896
rect 120718 239884 120724 239896
rect 117096 239856 120724 239884
rect 117096 239844 117102 239856
rect 120718 239844 120724 239856
rect 120776 239844 120782 239896
rect 179414 239844 179420 239896
rect 179472 239884 179478 239896
rect 301222 239884 301228 239896
rect 179472 239856 301228 239884
rect 179472 239844 179478 239856
rect 301222 239844 301228 239856
rect 301280 239844 301286 239896
rect 160738 239368 160744 239420
rect 160796 239408 160802 239420
rect 168006 239408 168012 239420
rect 160796 239380 168012 239408
rect 160796 239368 160802 239380
rect 168006 239368 168012 239380
rect 168064 239368 168070 239420
rect 310422 239368 310428 239420
rect 310480 239408 310486 239420
rect 331306 239408 331312 239420
rect 310480 239380 331312 239408
rect 310480 239368 310486 239380
rect 331306 239368 331312 239380
rect 331364 239368 331370 239420
rect 96430 239232 96436 239284
rect 96488 239272 96494 239284
rect 97718 239272 97724 239284
rect 96488 239244 97724 239272
rect 96488 239232 96494 239244
rect 97718 239232 97724 239244
rect 97776 239232 97782 239284
rect 82906 239096 82912 239148
rect 82964 239136 82970 239148
rect 292666 239136 292672 239148
rect 82964 239108 292672 239136
rect 82964 239096 82970 239108
rect 292666 239096 292672 239108
rect 292724 239096 292730 239148
rect 25498 239028 25504 239080
rect 25556 239068 25562 239080
rect 81434 239068 81440 239080
rect 25556 239040 81440 239068
rect 25556 239028 25562 239040
rect 81434 239028 81440 239040
rect 81492 239068 81498 239080
rect 82262 239068 82268 239080
rect 81492 239040 82268 239068
rect 81492 239028 81498 239040
rect 82262 239028 82268 239040
rect 82320 239028 82326 239080
rect 63494 238960 63500 239012
rect 63552 239000 63558 239012
rect 70026 239000 70032 239012
rect 63552 238972 70032 239000
rect 63552 238960 63558 238972
rect 70026 238960 70032 238972
rect 70084 238960 70090 239012
rect 107378 238960 107384 239012
rect 107436 239000 107442 239012
rect 139486 239000 139492 239012
rect 107436 238972 139492 239000
rect 107436 238960 107442 238972
rect 139486 238960 139492 238972
rect 139544 238960 139550 239012
rect 48130 238892 48136 238944
rect 48188 238932 48194 238944
rect 78674 238932 78680 238944
rect 48188 238904 78680 238932
rect 48188 238892 48194 238904
rect 78674 238892 78680 238904
rect 78732 238932 78738 238944
rect 79686 238932 79692 238944
rect 78732 238904 79692 238932
rect 78732 238892 78738 238904
rect 79686 238892 79692 238904
rect 79744 238892 79750 238944
rect 99374 238892 99380 238944
rect 99432 238932 99438 238944
rect 99650 238932 99656 238944
rect 99432 238904 99656 238932
rect 99432 238892 99438 238904
rect 99650 238892 99656 238904
rect 99708 238932 99714 238944
rect 135898 238932 135904 238944
rect 99708 238904 135904 238932
rect 99708 238892 99714 238904
rect 135898 238892 135904 238904
rect 135956 238892 135962 238944
rect 59078 238824 59084 238876
rect 59136 238864 59142 238876
rect 253014 238864 253020 238876
rect 59136 238836 253020 238864
rect 59136 238824 59142 238836
rect 253014 238824 253020 238836
rect 253072 238864 253078 238876
rect 298186 238864 298192 238876
rect 253072 238836 298192 238864
rect 253072 238824 253078 238836
rect 298186 238824 298192 238836
rect 298244 238824 298250 238876
rect 42518 238688 42524 238740
rect 42576 238728 42582 238740
rect 82906 238728 82912 238740
rect 42576 238700 82912 238728
rect 42576 238688 42582 238700
rect 82906 238688 82912 238700
rect 82964 238688 82970 238740
rect 119798 238688 119804 238740
rect 119856 238728 119862 238740
rect 124858 238728 124864 238740
rect 119856 238700 124864 238728
rect 119856 238688 119862 238700
rect 124858 238688 124864 238700
rect 124916 238688 124922 238740
rect 127526 238688 127532 238740
rect 127584 238728 127590 238740
rect 250530 238728 250536 238740
rect 127584 238700 250536 238728
rect 127584 238688 127590 238700
rect 250530 238688 250536 238700
rect 250588 238688 250594 238740
rect 265526 238688 265532 238740
rect 265584 238728 265590 238740
rect 299566 238728 299572 238740
rect 265584 238700 299572 238728
rect 265584 238688 265590 238700
rect 299566 238688 299572 238700
rect 299624 238688 299630 238740
rect 55122 238620 55128 238672
rect 55180 238660 55186 238672
rect 89346 238660 89352 238672
rect 55180 238632 89352 238660
rect 55180 238620 55186 238632
rect 89346 238620 89352 238632
rect 89404 238620 89410 238672
rect 91922 238620 91928 238672
rect 91980 238660 91986 238672
rect 149698 238660 149704 238672
rect 91980 238632 149704 238660
rect 91980 238620 91986 238632
rect 149698 238620 149704 238632
rect 149756 238620 149762 238672
rect 162302 238620 162308 238672
rect 162360 238660 162366 238672
rect 276014 238660 276020 238672
rect 162360 238632 276020 238660
rect 162360 238620 162366 238632
rect 276014 238620 276020 238632
rect 276072 238660 276078 238672
rect 310606 238660 310612 238672
rect 276072 238632 310612 238660
rect 276072 238620 276078 238632
rect 310606 238620 310612 238632
rect 310664 238620 310670 238672
rect 59170 238552 59176 238604
rect 59228 238592 59234 238604
rect 91278 238592 91284 238604
rect 59228 238564 91284 238592
rect 59228 238552 59234 238564
rect 91278 238552 91284 238564
rect 91336 238552 91342 238604
rect 105446 238552 105452 238604
rect 105504 238592 105510 238604
rect 173802 238592 173808 238604
rect 105504 238564 173808 238592
rect 105504 238552 105510 238564
rect 173802 238552 173808 238564
rect 173860 238552 173866 238604
rect 176010 238552 176016 238604
rect 176068 238592 176074 238604
rect 254394 238592 254400 238604
rect 176068 238564 254400 238592
rect 176068 238552 176074 238564
rect 254394 238552 254400 238564
rect 254452 238552 254458 238604
rect 288158 238552 288164 238604
rect 288216 238592 288222 238604
rect 313274 238592 313280 238604
rect 288216 238564 313280 238592
rect 288216 238552 288222 238564
rect 313274 238552 313280 238564
rect 313332 238552 313338 238604
rect 99006 238484 99012 238536
rect 99064 238524 99070 238536
rect 120902 238524 120908 238536
rect 99064 238496 120908 238524
rect 99064 238484 99070 238496
rect 120902 238484 120908 238496
rect 120960 238484 120966 238536
rect 169294 238484 169300 238536
rect 169352 238524 169358 238536
rect 204898 238524 204904 238536
rect 169352 238496 204904 238524
rect 169352 238484 169358 238496
rect 204898 238484 204904 238496
rect 204956 238484 204962 238536
rect 240778 238484 240784 238536
rect 240836 238524 240842 238536
rect 296070 238524 296076 238536
rect 240836 238496 296076 238524
rect 240836 238484 240842 238496
rect 296070 238484 296076 238496
rect 296128 238484 296134 238536
rect 117682 238416 117688 238468
rect 117740 238456 117746 238468
rect 127526 238456 127532 238468
rect 117740 238428 127532 238456
rect 117740 238416 117746 238428
rect 127526 238416 127532 238428
rect 127584 238416 127590 238468
rect 174630 238416 174636 238468
rect 174688 238456 174694 238468
rect 195974 238456 195980 238468
rect 174688 238428 195980 238456
rect 174688 238416 174694 238428
rect 195974 238416 195980 238428
rect 196032 238416 196038 238468
rect 88058 238348 88064 238400
rect 88116 238388 88122 238400
rect 91738 238388 91744 238400
rect 88116 238360 91744 238388
rect 88116 238348 88122 238360
rect 91738 238348 91744 238360
rect 91796 238348 91802 238400
rect 108942 238348 108948 238400
rect 109000 238388 109006 238400
rect 123478 238388 123484 238400
rect 109000 238360 123484 238388
rect 109000 238348 109006 238360
rect 123478 238348 123484 238360
rect 123536 238348 123542 238400
rect 96522 238280 96528 238332
rect 96580 238320 96586 238332
rect 119890 238320 119896 238332
rect 96580 238292 119896 238320
rect 96580 238280 96586 238292
rect 119890 238280 119896 238292
rect 119948 238280 119954 238332
rect 60642 238144 60648 238196
rect 60700 238184 60706 238196
rect 73062 238184 73068 238196
rect 60700 238156 73068 238184
rect 60700 238144 60706 238156
rect 73062 238144 73068 238156
rect 73120 238184 73126 238196
rect 73890 238184 73896 238196
rect 73120 238156 73896 238184
rect 73120 238144 73126 238156
rect 73890 238144 73896 238156
rect 73948 238144 73954 238196
rect 71314 238076 71320 238128
rect 71372 238116 71378 238128
rect 86218 238116 86224 238128
rect 71372 238088 86224 238116
rect 71372 238076 71378 238088
rect 86218 238076 86224 238088
rect 86276 238076 86282 238128
rect 93210 238076 93216 238128
rect 93268 238116 93274 238128
rect 98822 238116 98828 238128
rect 93268 238088 98828 238116
rect 93268 238076 93274 238088
rect 98822 238076 98828 238088
rect 98880 238076 98886 238128
rect 195974 238076 195980 238128
rect 196032 238116 196038 238128
rect 210602 238116 210608 238128
rect 196032 238088 210608 238116
rect 196032 238076 196038 238088
rect 210602 238076 210608 238088
rect 210660 238076 210666 238128
rect 57882 238008 57888 238060
rect 57940 238048 57946 238060
rect 92474 238048 92480 238060
rect 57940 238020 92480 238048
rect 57940 238008 57946 238020
rect 92474 238008 92480 238020
rect 92532 238008 92538 238060
rect 122282 238008 122288 238060
rect 122340 238048 122346 238060
rect 327166 238048 327172 238060
rect 122340 238020 327172 238048
rect 122340 238008 122346 238020
rect 327166 238008 327172 238020
rect 327224 238008 327230 238060
rect 108022 237940 108028 237992
rect 108080 237980 108086 237992
rect 108942 237980 108948 237992
rect 108080 237952 108948 237980
rect 108080 237940 108086 237952
rect 108942 237940 108948 237952
rect 109000 237940 109006 237992
rect 92474 237464 92480 237516
rect 92532 237504 92538 237516
rect 93762 237504 93768 237516
rect 92532 237476 93768 237504
rect 92532 237464 92538 237476
rect 93762 237464 93768 237476
rect 93820 237504 93826 237516
rect 95142 237504 95148 237516
rect 93820 237476 95148 237504
rect 93820 237464 93826 237476
rect 95142 237464 95148 237476
rect 95200 237464 95206 237516
rect 70026 237396 70032 237448
rect 70084 237436 70090 237448
rect 71038 237436 71044 237448
rect 70084 237408 71044 237436
rect 70084 237396 70090 237408
rect 71038 237396 71044 237408
rect 71096 237396 71102 237448
rect 75546 237396 75552 237448
rect 75604 237436 75610 237448
rect 77110 237436 77116 237448
rect 75604 237408 77116 237436
rect 75604 237396 75610 237408
rect 77110 237396 77116 237408
rect 77168 237396 77174 237448
rect 103514 237436 103520 237448
rect 93826 237408 103520 237436
rect 2958 237328 2964 237380
rect 3016 237368 3022 237380
rect 93826 237368 93854 237408
rect 103514 237396 103520 237408
rect 103572 237436 103578 237448
rect 104526 237436 104532 237448
rect 103572 237408 104532 237436
rect 103572 237396 103578 237408
rect 104526 237396 104532 237408
rect 104584 237396 104590 237448
rect 104618 237396 104624 237448
rect 104676 237436 104682 237448
rect 106090 237436 106096 237448
rect 104676 237408 106096 237436
rect 104676 237396 104682 237408
rect 106090 237396 106096 237408
rect 106148 237396 106154 237448
rect 173802 237396 173808 237448
rect 173860 237436 173866 237448
rect 175918 237436 175924 237448
rect 173860 237408 175924 237436
rect 173860 237396 173866 237408
rect 175918 237396 175924 237408
rect 175976 237396 175982 237448
rect 209314 237396 209320 237448
rect 209372 237436 209378 237448
rect 210418 237436 210424 237448
rect 209372 237408 210424 237436
rect 209372 237396 209378 237408
rect 210418 237396 210424 237408
rect 210476 237396 210482 237448
rect 213178 237396 213184 237448
rect 213236 237436 213242 237448
rect 216030 237436 216036 237448
rect 213236 237408 216036 237436
rect 213236 237396 213242 237408
rect 216030 237396 216036 237408
rect 216088 237396 216094 237448
rect 265618 237396 265624 237448
rect 265676 237436 265682 237448
rect 267274 237436 267280 237448
rect 265676 237408 267280 237436
rect 265676 237396 265682 237408
rect 267274 237396 267280 237408
rect 267332 237396 267338 237448
rect 283558 237396 283564 237448
rect 283616 237436 283622 237448
rect 284294 237436 284300 237448
rect 283616 237408 284300 237436
rect 283616 237396 283622 237408
rect 284294 237396 284300 237408
rect 284352 237396 284358 237448
rect 291930 237396 291936 237448
rect 291988 237436 291994 237448
rect 292574 237436 292580 237448
rect 291988 237408 292580 237436
rect 291988 237396 291994 237408
rect 292574 237396 292580 237408
rect 292632 237396 292638 237448
rect 3016 237340 93854 237368
rect 3016 237328 3022 237340
rect 122466 237328 122472 237380
rect 122524 237368 122530 237380
rect 322934 237368 322940 237380
rect 122524 237340 322940 237368
rect 122524 237328 122530 237340
rect 322934 237328 322940 237340
rect 322992 237328 322998 237380
rect 46658 237260 46664 237312
rect 46716 237300 46722 237312
rect 106734 237300 106740 237312
rect 46716 237272 106740 237300
rect 46716 237260 46722 237272
rect 106734 237260 106740 237272
rect 106792 237300 106798 237312
rect 123570 237300 123576 237312
rect 106792 237272 123576 237300
rect 106792 237260 106798 237272
rect 123570 237260 123576 237272
rect 123628 237260 123634 237312
rect 145650 237260 145656 237312
rect 145708 237300 145714 237312
rect 296898 237300 296904 237312
rect 145708 237272 296904 237300
rect 145708 237260 145714 237272
rect 296898 237260 296904 237272
rect 296956 237260 296962 237312
rect 45370 237192 45376 237244
rect 45428 237232 45434 237244
rect 81618 237232 81624 237244
rect 45428 237204 81624 237232
rect 45428 237192 45434 237204
rect 81618 237192 81624 237204
rect 81676 237192 81682 237244
rect 95786 237192 95792 237244
rect 95844 237232 95850 237244
rect 152458 237232 152464 237244
rect 95844 237204 152464 237232
rect 95844 237192 95850 237204
rect 152458 237192 152464 237204
rect 152516 237192 152522 237244
rect 162394 237192 162400 237244
rect 162452 237232 162458 237244
rect 302418 237232 302424 237244
rect 162452 237204 302424 237232
rect 162452 237192 162458 237204
rect 302418 237192 302424 237204
rect 302476 237192 302482 237244
rect 41138 237124 41144 237176
rect 41196 237164 41202 237176
rect 73246 237164 73252 237176
rect 41196 237136 73252 237164
rect 41196 237124 41202 237136
rect 73246 237124 73252 237136
rect 73304 237124 73310 237176
rect 98822 237124 98828 237176
rect 98880 237164 98886 237176
rect 99282 237164 99288 237176
rect 98880 237136 99288 237164
rect 98880 237124 98886 237136
rect 99282 237124 99288 237136
rect 99340 237164 99346 237176
rect 126422 237164 126428 237176
rect 99340 237136 126428 237164
rect 99340 237124 99346 237136
rect 126422 237124 126428 237136
rect 126480 237124 126486 237176
rect 159358 237124 159364 237176
rect 159416 237164 159422 237176
rect 269206 237164 269212 237176
rect 159416 237136 269212 237164
rect 159416 237124 159422 237136
rect 269206 237124 269212 237136
rect 269264 237124 269270 237176
rect 290458 237124 290464 237176
rect 290516 237164 290522 237176
rect 300854 237164 300860 237176
rect 290516 237136 300860 237164
rect 290516 237124 290522 237136
rect 300854 237124 300860 237136
rect 300912 237124 300918 237176
rect 158162 237056 158168 237108
rect 158220 237096 158226 237108
rect 191926 237096 191932 237108
rect 158220 237068 191932 237096
rect 158220 237056 158226 237068
rect 191926 237056 191932 237068
rect 191984 237056 191990 237108
rect 233878 237056 233884 237108
rect 233936 237096 233942 237108
rect 299474 237096 299480 237108
rect 233936 237068 299480 237096
rect 233936 237056 233942 237068
rect 299474 237056 299480 237068
rect 299532 237056 299538 237108
rect 141510 236648 141516 236700
rect 141568 236688 141574 236700
rect 239490 236688 239496 236700
rect 141568 236660 239496 236688
rect 141568 236648 141574 236660
rect 239490 236648 239496 236660
rect 239548 236648 239554 236700
rect 278774 236648 278780 236700
rect 278832 236688 278838 236700
rect 294230 236688 294236 236700
rect 278832 236660 294236 236688
rect 278832 236648 278838 236660
rect 294230 236648 294236 236660
rect 294288 236648 294294 236700
rect 73246 235968 73252 236020
rect 73304 236008 73310 236020
rect 73798 236008 73804 236020
rect 73304 235980 73804 236008
rect 73304 235968 73310 235980
rect 73798 235968 73804 235980
rect 73856 235968 73862 236020
rect 322934 235968 322940 236020
rect 322992 236008 322998 236020
rect 323578 236008 323584 236020
rect 322992 235980 323584 236008
rect 322992 235968 322998 235980
rect 323578 235968 323584 235980
rect 323636 235968 323642 236020
rect 46750 235900 46756 235952
rect 46808 235940 46814 235952
rect 302326 235940 302332 235952
rect 46808 235912 302332 235940
rect 46808 235900 46814 235912
rect 302326 235900 302332 235912
rect 302384 235900 302390 235952
rect 26878 235832 26884 235884
rect 26936 235872 26942 235884
rect 112530 235872 112536 235884
rect 26936 235844 112536 235872
rect 26936 235832 26942 235844
rect 112530 235832 112536 235844
rect 112588 235872 112594 235884
rect 131114 235872 131120 235884
rect 112588 235844 131120 235872
rect 112588 235832 112594 235844
rect 131114 235832 131120 235844
rect 131172 235832 131178 235884
rect 176102 235832 176108 235884
rect 176160 235872 176166 235884
rect 274082 235872 274088 235884
rect 176160 235844 274088 235872
rect 176160 235832 176166 235844
rect 274082 235832 274088 235844
rect 274140 235872 274146 235884
rect 306466 235872 306472 235884
rect 274140 235844 306472 235872
rect 274140 235832 274146 235844
rect 306466 235832 306472 235844
rect 306524 235832 306530 235884
rect 52362 235764 52368 235816
rect 52420 235804 52426 235816
rect 80330 235804 80336 235816
rect 52420 235776 80336 235804
rect 52420 235764 52426 235776
rect 80330 235764 80336 235776
rect 80388 235764 80394 235816
rect 88242 235764 88248 235816
rect 88300 235804 88306 235816
rect 126974 235804 126980 235816
rect 88300 235776 126980 235804
rect 88300 235764 88306 235776
rect 126974 235764 126980 235776
rect 127032 235764 127038 235816
rect 46842 235696 46848 235748
rect 46900 235736 46906 235748
rect 71958 235736 71964 235748
rect 46900 235708 71964 235736
rect 46900 235696 46906 235708
rect 71958 235696 71964 235708
rect 72016 235696 72022 235748
rect 87414 235356 87420 235408
rect 87472 235396 87478 235408
rect 88242 235396 88248 235408
rect 87472 235368 88248 235396
rect 87472 235356 87478 235368
rect 88242 235356 88248 235368
rect 88300 235356 88306 235408
rect 129642 235396 129648 235408
rect 122806 235368 129648 235396
rect 102226 235288 102232 235340
rect 102284 235328 102290 235340
rect 122806 235328 122834 235368
rect 129642 235356 129648 235368
rect 129700 235396 129706 235408
rect 130562 235396 130568 235408
rect 129700 235368 130568 235396
rect 129700 235356 129706 235368
rect 130562 235356 130568 235368
rect 130620 235356 130626 235408
rect 166718 235356 166724 235408
rect 166776 235396 166782 235408
rect 192478 235396 192484 235408
rect 166776 235368 192484 235396
rect 166776 235356 166782 235368
rect 192478 235356 192484 235368
rect 192536 235356 192542 235408
rect 102284 235300 122834 235328
rect 102284 235288 102290 235300
rect 151262 235288 151268 235340
rect 151320 235328 151326 235340
rect 244918 235328 244924 235340
rect 151320 235300 244924 235328
rect 151320 235288 151326 235300
rect 244918 235288 244924 235300
rect 244976 235288 244982 235340
rect 60550 235220 60556 235272
rect 60608 235260 60614 235272
rect 247678 235260 247684 235272
rect 60608 235232 247684 235260
rect 60608 235220 60614 235232
rect 247678 235220 247684 235232
rect 247736 235220 247742 235272
rect 250530 235220 250536 235272
rect 250588 235260 250594 235272
rect 353938 235260 353944 235272
rect 250588 235232 353944 235260
rect 250588 235220 250594 235232
rect 353938 235220 353944 235232
rect 353996 235220 354002 235272
rect 46198 234608 46204 234660
rect 46256 234648 46262 234660
rect 46750 234648 46756 234660
rect 46256 234620 46756 234648
rect 46256 234608 46262 234620
rect 46750 234608 46756 234620
rect 46808 234608 46814 234660
rect 71958 234608 71964 234660
rect 72016 234648 72022 234660
rect 72418 234648 72424 234660
rect 72016 234620 72424 234648
rect 72016 234608 72022 234620
rect 72418 234608 72424 234620
rect 72476 234608 72482 234660
rect 80330 234608 80336 234660
rect 80388 234648 80394 234660
rect 80698 234648 80704 234660
rect 80388 234620 80704 234648
rect 80388 234608 80394 234620
rect 80698 234608 80704 234620
rect 80756 234608 80762 234660
rect 56318 234540 56324 234592
rect 56376 234580 56382 234592
rect 349246 234580 349252 234592
rect 56376 234552 349252 234580
rect 56376 234540 56382 234552
rect 349246 234540 349252 234552
rect 349304 234540 349310 234592
rect 63402 234472 63408 234524
rect 63460 234512 63466 234524
rect 265526 234512 265532 234524
rect 63460 234484 265532 234512
rect 63460 234472 63466 234484
rect 265526 234472 265532 234484
rect 265584 234472 265590 234524
rect 317414 234512 317420 234524
rect 296686 234484 317420 234512
rect 13078 234404 13084 234456
rect 13136 234444 13142 234456
rect 86862 234444 86868 234456
rect 13136 234416 86868 234444
rect 13136 234404 13142 234416
rect 86862 234404 86868 234416
rect 86920 234404 86926 234456
rect 110598 234404 110604 234456
rect 110656 234444 110662 234456
rect 111058 234444 111064 234456
rect 110656 234416 111064 234444
rect 110656 234404 110662 234416
rect 111058 234404 111064 234416
rect 111116 234444 111122 234456
rect 129090 234444 129096 234456
rect 111116 234416 129096 234444
rect 111116 234404 111122 234416
rect 129090 234404 129096 234416
rect 129148 234404 129154 234456
rect 166350 234404 166356 234456
rect 166408 234444 166414 234456
rect 296686 234444 296714 234484
rect 317414 234472 317420 234484
rect 317472 234512 317478 234524
rect 318058 234512 318064 234524
rect 317472 234484 318064 234512
rect 317472 234472 317478 234484
rect 318058 234472 318064 234484
rect 318116 234472 318122 234524
rect 166408 234416 296714 234444
rect 166408 234404 166414 234416
rect 83458 234336 83464 234388
rect 83516 234376 83522 234388
rect 144178 234376 144184 234388
rect 83516 234348 144184 234376
rect 83516 234336 83522 234348
rect 144178 234336 144184 234348
rect 144236 234336 144242 234388
rect 160922 233996 160928 234048
rect 160980 234036 160986 234048
rect 214558 234036 214564 234048
rect 160980 234008 214564 234036
rect 160980 233996 160986 234008
rect 214558 233996 214564 234008
rect 214616 233996 214622 234048
rect 171962 233928 171968 233980
rect 172020 233968 172026 233980
rect 264330 233968 264336 233980
rect 172020 233940 264336 233968
rect 172020 233928 172026 233940
rect 264330 233928 264336 233940
rect 264388 233928 264394 233980
rect 84194 233860 84200 233912
rect 84252 233900 84258 233912
rect 84838 233900 84844 233912
rect 84252 233872 84844 233900
rect 84252 233860 84258 233872
rect 84838 233860 84844 233872
rect 84896 233860 84902 233912
rect 89714 233860 89720 233912
rect 89772 233900 89778 233912
rect 90634 233900 90640 233912
rect 89772 233872 90640 233900
rect 89772 233860 89778 233872
rect 90634 233860 90640 233872
rect 90692 233860 90698 233912
rect 93946 233860 93952 233912
rect 94004 233900 94010 233912
rect 94498 233900 94504 233912
rect 94004 233872 94504 233900
rect 94004 233860 94010 233872
rect 94498 233860 94504 233872
rect 94556 233860 94562 233912
rect 100754 233860 100760 233912
rect 100812 233900 100818 233912
rect 101582 233900 101588 233912
rect 100812 233872 101588 233900
rect 100812 233860 100818 233872
rect 101582 233860 101588 233872
rect 101640 233860 101646 233912
rect 103698 233860 103704 233912
rect 103756 233900 103762 233912
rect 104802 233900 104808 233912
rect 103756 233872 104808 233900
rect 103756 233860 103762 233872
rect 104802 233860 104808 233872
rect 104860 233860 104866 233912
rect 114554 233860 114560 233912
rect 114612 233900 114618 233912
rect 115750 233900 115756 233912
rect 114612 233872 115756 233900
rect 114612 233860 114618 233872
rect 115750 233860 115756 233872
rect 115808 233860 115814 233912
rect 169202 233860 169208 233912
rect 169260 233900 169266 233912
rect 324590 233900 324596 233912
rect 169260 233872 324596 233900
rect 169260 233860 169266 233872
rect 324590 233860 324596 233872
rect 324648 233860 324654 233912
rect 114462 233248 114468 233300
rect 114520 233288 114526 233300
rect 117958 233288 117964 233300
rect 114520 233260 117964 233288
rect 114520 233248 114526 233260
rect 117958 233248 117964 233260
rect 118016 233248 118022 233300
rect 61838 233180 61844 233232
rect 61896 233220 61902 233232
rect 288158 233220 288164 233232
rect 61896 233192 288164 233220
rect 61896 233180 61902 233192
rect 288158 233180 288164 233192
rect 288216 233180 288222 233232
rect 347038 233180 347044 233232
rect 347096 233220 347102 233232
rect 580166 233220 580172 233232
rect 347096 233192 580172 233220
rect 347096 233180 347102 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 113818 233112 113824 233164
rect 113876 233152 113882 233164
rect 296806 233152 296812 233164
rect 113876 233124 296812 233152
rect 113876 233112 113882 233124
rect 296806 233112 296812 233124
rect 296864 233112 296870 233164
rect 45278 233044 45284 233096
rect 45336 233084 45342 233096
rect 75178 233084 75184 233096
rect 45336 233056 75184 233084
rect 45336 233044 45342 233056
rect 75178 233044 75184 233056
rect 75236 233084 75242 233096
rect 75546 233084 75552 233096
rect 75236 233056 75552 233084
rect 75236 233044 75242 233056
rect 75546 233044 75552 233056
rect 75604 233044 75610 233096
rect 76466 233044 76472 233096
rect 76524 233084 76530 233096
rect 137278 233084 137284 233096
rect 76524 233056 137284 233084
rect 76524 233044 76530 233056
rect 137278 233044 137284 233056
rect 137336 233044 137342 233096
rect 148594 233044 148600 233096
rect 148652 233084 148658 233096
rect 295518 233084 295524 233096
rect 148652 233056 295524 233084
rect 148652 233044 148658 233056
rect 295518 233044 295524 233056
rect 295576 233044 295582 233096
rect 44082 232976 44088 233028
rect 44140 233016 44146 233028
rect 77754 233016 77760 233028
rect 44140 232988 77760 233016
rect 44140 232976 44146 232988
rect 77754 232976 77760 232988
rect 77812 233016 77818 233028
rect 77938 233016 77944 233028
rect 77812 232988 77944 233016
rect 77812 232976 77818 232988
rect 77938 232976 77944 232988
rect 77996 232976 78002 233028
rect 86862 232976 86868 233028
rect 86920 233016 86926 233028
rect 195974 233016 195980 233028
rect 86920 232988 195980 233016
rect 86920 232976 86926 232988
rect 195974 232976 195980 232988
rect 196032 232976 196038 233028
rect 27522 232908 27528 232960
rect 27580 232948 27586 232960
rect 113174 232948 113180 232960
rect 27580 232920 113180 232948
rect 27580 232908 27586 232920
rect 113174 232908 113180 232920
rect 113232 232948 113238 232960
rect 114462 232948 114468 232960
rect 113232 232920 114468 232948
rect 113232 232908 113238 232920
rect 114462 232908 114468 232920
rect 114520 232908 114526 232960
rect 167914 232908 167920 232960
rect 167972 232948 167978 232960
rect 271138 232948 271144 232960
rect 167972 232920 271144 232948
rect 167972 232908 167978 232920
rect 271138 232908 271144 232920
rect 271196 232908 271202 232960
rect 311158 232568 311164 232620
rect 311216 232608 311222 232620
rect 335446 232608 335452 232620
rect 311216 232580 335452 232608
rect 311216 232568 311222 232580
rect 335446 232568 335452 232580
rect 335504 232568 335510 232620
rect 282178 232500 282184 232552
rect 282236 232540 282242 232552
rect 313366 232540 313372 232552
rect 282236 232512 313372 232540
rect 282236 232500 282242 232512
rect 313366 232500 313372 232512
rect 313424 232500 313430 232552
rect 128354 231820 128360 231872
rect 128412 231860 128418 231872
rect 128998 231860 129004 231872
rect 128412 231832 129004 231860
rect 128412 231820 128418 231832
rect 128998 231820 129004 231832
rect 129056 231860 129062 231872
rect 346578 231860 346584 231872
rect 129056 231832 346584 231860
rect 129056 231820 129062 231832
rect 346578 231820 346584 231832
rect 346636 231820 346642 231872
rect 61930 231752 61936 231804
rect 61988 231792 61994 231804
rect 298370 231792 298376 231804
rect 61988 231764 298376 231792
rect 61988 231752 61994 231764
rect 298370 231752 298376 231764
rect 298428 231752 298434 231804
rect 81618 231684 81624 231736
rect 81676 231724 81682 231736
rect 278866 231724 278872 231736
rect 81676 231696 278872 231724
rect 81676 231684 81682 231696
rect 278866 231684 278872 231696
rect 278924 231684 278930 231736
rect 37090 231616 37096 231668
rect 37148 231656 37154 231668
rect 104250 231656 104256 231668
rect 37148 231628 104256 231656
rect 37148 231616 37154 231628
rect 104250 231616 104256 231628
rect 104308 231656 104314 231668
rect 104618 231656 104624 231668
rect 104308 231628 104624 231656
rect 104308 231616 104314 231628
rect 104618 231616 104624 231628
rect 104676 231616 104682 231668
rect 169754 231616 169760 231668
rect 169812 231656 169818 231668
rect 171042 231656 171048 231668
rect 169812 231628 171048 231656
rect 169812 231616 169818 231628
rect 171042 231616 171048 231628
rect 171100 231656 171106 231668
rect 305270 231656 305276 231668
rect 171100 231628 305276 231656
rect 171100 231616 171106 231628
rect 305270 231616 305276 231628
rect 305328 231616 305334 231668
rect 115106 231548 115112 231600
rect 115164 231588 115170 231600
rect 179782 231588 179788 231600
rect 115164 231560 179788 231588
rect 115164 231548 115170 231560
rect 179782 231548 179788 231560
rect 179840 231588 179846 231600
rect 235994 231588 236000 231600
rect 179840 231560 236000 231588
rect 179840 231548 179846 231560
rect 235994 231548 236000 231560
rect 236052 231548 236058 231600
rect 88702 231480 88708 231532
rect 88760 231520 88766 231532
rect 128354 231520 128360 231532
rect 88760 231492 128360 231520
rect 88760 231480 88766 231492
rect 128354 231480 128360 231492
rect 128412 231480 128418 231532
rect 154482 231140 154488 231192
rect 154540 231180 154546 231192
rect 169754 231180 169760 231192
rect 154540 231152 169760 231180
rect 154540 231140 154546 231152
rect 169754 231140 169760 231152
rect 169812 231140 169818 231192
rect 173250 231140 173256 231192
rect 173308 231180 173314 231192
rect 222838 231180 222844 231192
rect 173308 231152 222844 231180
rect 173308 231140 173314 231152
rect 222838 231140 222844 231152
rect 222896 231140 222902 231192
rect 68738 231072 68744 231124
rect 68796 231112 68802 231124
rect 325786 231112 325792 231124
rect 68796 231084 325792 231112
rect 68796 231072 68802 231084
rect 325786 231072 325792 231084
rect 325844 231072 325850 231124
rect 39758 230392 39764 230444
rect 39816 230432 39822 230444
rect 104158 230432 104164 230444
rect 39816 230404 104164 230432
rect 39816 230392 39822 230404
rect 104158 230392 104164 230404
rect 104216 230392 104222 230444
rect 104526 230392 104532 230444
rect 104584 230432 104590 230444
rect 154482 230432 154488 230444
rect 104584 230404 154488 230432
rect 104584 230392 104590 230404
rect 154482 230392 154488 230404
rect 154540 230392 154546 230444
rect 172054 230392 172060 230444
rect 172112 230432 172118 230444
rect 332594 230432 332600 230444
rect 172112 230404 332600 230432
rect 172112 230392 172118 230404
rect 332594 230392 332600 230404
rect 332652 230392 332658 230444
rect 98362 230324 98368 230376
rect 98420 230364 98426 230376
rect 233878 230364 233884 230376
rect 98420 230336 233884 230364
rect 98420 230324 98426 230336
rect 233878 230324 233884 230336
rect 233936 230324 233942 230376
rect 118326 230256 118332 230308
rect 118384 230296 118390 230308
rect 240778 230296 240784 230308
rect 118384 230268 240784 230296
rect 118384 230256 118390 230268
rect 240778 230256 240784 230268
rect 240836 230256 240842 230308
rect 63218 229780 63224 229832
rect 63276 229820 63282 229832
rect 161474 229820 161480 229832
rect 63276 229792 161480 229820
rect 63276 229780 63282 229792
rect 161474 229780 161480 229792
rect 161532 229780 161538 229832
rect 161382 229712 161388 229764
rect 161440 229752 161446 229764
rect 574738 229752 574744 229764
rect 161440 229724 574744 229752
rect 161440 229712 161446 229724
rect 574738 229712 574744 229724
rect 574796 229712 574802 229764
rect 74718 229032 74724 229084
rect 74776 229072 74782 229084
rect 294138 229072 294144 229084
rect 74776 229044 294144 229072
rect 74776 229032 74782 229044
rect 294138 229032 294144 229044
rect 294196 229032 294202 229084
rect 38562 228964 38568 229016
rect 38620 229004 38626 229016
rect 122926 229004 122932 229016
rect 38620 228976 122932 229004
rect 38620 228964 38626 228976
rect 122926 228964 122932 228976
rect 122984 228964 122990 229016
rect 155218 228964 155224 229016
rect 155276 229004 155282 229016
rect 328546 229004 328552 229016
rect 155276 228976 328552 229004
rect 155276 228964 155282 228976
rect 328546 228964 328552 228976
rect 328604 228964 328610 229016
rect 69106 228896 69112 228948
rect 69164 228936 69170 228948
rect 241514 228936 241520 228948
rect 69164 228908 241520 228936
rect 69164 228896 69170 228908
rect 241514 228896 241520 228908
rect 241572 228896 241578 228948
rect 159450 228352 159456 228404
rect 159508 228392 159514 228404
rect 255314 228392 255320 228404
rect 159508 228364 255320 228392
rect 159508 228352 159514 228364
rect 255314 228352 255320 228364
rect 255372 228352 255378 228404
rect 122926 227740 122932 227792
rect 122984 227780 122990 227792
rect 124858 227780 124864 227792
rect 122984 227752 124864 227780
rect 122984 227740 122990 227752
rect 124858 227740 124864 227752
rect 124916 227740 124922 227792
rect 53650 227672 53656 227724
rect 53708 227712 53714 227724
rect 287698 227712 287704 227724
rect 53708 227684 287704 227712
rect 53708 227672 53714 227684
rect 287698 227672 287704 227684
rect 287756 227672 287762 227724
rect 108666 227604 108672 227656
rect 108724 227644 108730 227656
rect 153102 227644 153108 227656
rect 108724 227616 153108 227644
rect 108724 227604 108730 227616
rect 153102 227604 153108 227616
rect 153160 227604 153166 227656
rect 163498 227604 163504 227656
rect 163556 227644 163562 227656
rect 218054 227644 218060 227656
rect 163556 227616 218060 227644
rect 163556 227604 163562 227616
rect 218054 227604 218060 227616
rect 218112 227604 218118 227656
rect 145558 227196 145564 227248
rect 145616 227236 145622 227248
rect 232498 227236 232504 227248
rect 145616 227208 232504 227236
rect 145616 227196 145622 227208
rect 232498 227196 232504 227208
rect 232556 227196 232562 227248
rect 100938 227128 100944 227180
rect 100996 227168 101002 227180
rect 198182 227168 198188 227180
rect 100996 227140 198188 227168
rect 100996 227128 101002 227140
rect 198182 227128 198188 227140
rect 198240 227128 198246 227180
rect 60458 227060 60464 227112
rect 60516 227100 60522 227112
rect 158162 227100 158168 227112
rect 60516 227072 158168 227100
rect 60516 227060 60522 227072
rect 158162 227060 158168 227072
rect 158220 227060 158226 227112
rect 231854 227060 231860 227112
rect 231912 227100 231918 227112
rect 268378 227100 268384 227112
rect 231912 227072 268384 227100
rect 231912 227060 231918 227072
rect 268378 227060 268384 227072
rect 268436 227060 268442 227112
rect 153102 226992 153108 227044
rect 153160 227032 153166 227044
rect 329926 227032 329932 227044
rect 153160 227004 329932 227032
rect 153160 226992 153166 227004
rect 329926 226992 329932 227004
rect 329984 226992 329990 227044
rect 63310 226244 63316 226296
rect 63368 226284 63374 226296
rect 290458 226284 290464 226296
rect 63368 226256 290464 226284
rect 63368 226244 63374 226256
rect 290458 226244 290464 226256
rect 290516 226244 290522 226296
rect 177666 225632 177672 225684
rect 177724 225672 177730 225684
rect 189718 225672 189724 225684
rect 177724 225644 189724 225672
rect 177724 225632 177730 225644
rect 189718 225632 189724 225644
rect 189776 225632 189782 225684
rect 148318 225564 148324 225616
rect 148376 225604 148382 225616
rect 240778 225604 240784 225616
rect 148376 225576 240784 225604
rect 148376 225564 148382 225576
rect 240778 225564 240784 225576
rect 240836 225564 240842 225616
rect 325050 225564 325056 225616
rect 325108 225604 325114 225616
rect 332594 225604 332600 225616
rect 325108 225576 332600 225604
rect 325108 225564 325114 225576
rect 332594 225564 332600 225576
rect 332652 225564 332658 225616
rect 81434 224884 81440 224936
rect 81492 224924 81498 224936
rect 277394 224924 277400 224936
rect 81492 224896 277400 224924
rect 81492 224884 81498 224896
rect 277394 224884 277400 224896
rect 277452 224884 277458 224936
rect 3418 224204 3424 224256
rect 3476 224244 3482 224256
rect 120166 224244 120172 224256
rect 3476 224216 120172 224244
rect 3476 224204 3482 224216
rect 120166 224204 120172 224216
rect 120224 224204 120230 224256
rect 136174 224204 136180 224256
rect 136232 224244 136238 224256
rect 239398 224244 239404 224256
rect 136232 224216 239404 224244
rect 136232 224204 136238 224216
rect 239398 224204 239404 224216
rect 239456 224204 239462 224256
rect 68830 223524 68836 223576
rect 68888 223564 68894 223576
rect 324314 223564 324320 223576
rect 68888 223536 324320 223564
rect 68888 223524 68894 223536
rect 324314 223524 324320 223536
rect 324372 223524 324378 223576
rect 140222 222912 140228 222964
rect 140280 222952 140286 222964
rect 287790 222952 287796 222964
rect 140280 222924 287796 222952
rect 140280 222912 140286 222924
rect 287790 222912 287796 222924
rect 287848 222912 287854 222964
rect 79042 222844 79048 222896
rect 79100 222884 79106 222896
rect 273254 222884 273260 222896
rect 79100 222856 273260 222884
rect 79100 222844 79106 222856
rect 273254 222844 273260 222856
rect 273312 222844 273318 222896
rect 325142 222844 325148 222896
rect 325200 222884 325206 222896
rect 333974 222884 333980 222896
rect 325200 222856 333980 222884
rect 325200 222844 325206 222856
rect 333974 222844 333980 222856
rect 334032 222844 334038 222896
rect 170398 221484 170404 221536
rect 170456 221524 170462 221536
rect 203518 221524 203524 221536
rect 170456 221496 203524 221524
rect 170456 221484 170462 221496
rect 203518 221484 203524 221496
rect 203576 221484 203582 221536
rect 64598 221416 64604 221468
rect 64656 221456 64662 221468
rect 343634 221456 343640 221468
rect 64656 221428 343640 221456
rect 64656 221416 64662 221428
rect 343634 221416 343640 221428
rect 343692 221416 343698 221468
rect 58710 220192 58716 220244
rect 58768 220232 58774 220244
rect 122098 220232 122104 220244
rect 58768 220204 122104 220232
rect 58768 220192 58774 220204
rect 122098 220192 122104 220204
rect 122156 220192 122162 220244
rect 141602 220192 141608 220244
rect 141660 220232 141666 220244
rect 283650 220232 283656 220244
rect 141660 220204 283656 220232
rect 141660 220192 141666 220204
rect 283650 220192 283656 220204
rect 283708 220192 283714 220244
rect 89990 220124 89996 220176
rect 90048 220164 90054 220176
rect 252830 220164 252836 220176
rect 90048 220136 252836 220164
rect 90048 220124 90054 220136
rect 252830 220124 252836 220136
rect 252888 220124 252894 220176
rect 65978 220056 65984 220108
rect 66036 220096 66042 220108
rect 251174 220096 251180 220108
rect 66036 220068 251180 220096
rect 66036 220056 66042 220068
rect 251174 220056 251180 220068
rect 251232 220056 251238 220108
rect 256694 220056 256700 220108
rect 256752 220096 256758 220108
rect 278038 220096 278044 220108
rect 256752 220068 278044 220096
rect 256752 220056 256758 220068
rect 278038 220056 278044 220068
rect 278096 220056 278102 220108
rect 239490 219376 239496 219428
rect 239548 219416 239554 219428
rect 327074 219416 327080 219428
rect 239548 219388 327080 219416
rect 239548 219376 239554 219388
rect 327074 219376 327080 219388
rect 327132 219416 327138 219428
rect 335354 219416 335360 219428
rect 327132 219388 335360 219416
rect 327132 219376 327138 219388
rect 335354 219376 335360 219388
rect 335412 219376 335418 219428
rect 355318 219376 355324 219428
rect 355376 219416 355382 219428
rect 580166 219416 580172 219428
rect 355376 219388 580172 219416
rect 355376 219376 355382 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 52270 218900 52276 218952
rect 52328 218940 52334 218952
rect 163498 218940 163504 218952
rect 52328 218912 163504 218940
rect 52328 218900 52334 218912
rect 163498 218900 163504 218912
rect 163556 218900 163562 218952
rect 164970 218900 164976 218952
rect 165028 218940 165034 218952
rect 269114 218940 269120 218952
rect 165028 218912 269120 218940
rect 165028 218900 165034 218912
rect 269114 218900 269120 218912
rect 269172 218900 269178 218952
rect 99466 218832 99472 218884
rect 99524 218872 99530 218884
rect 220078 218872 220084 218884
rect 99524 218844 220084 218872
rect 99524 218832 99530 218844
rect 220078 218832 220084 218844
rect 220136 218832 220142 218884
rect 142890 218764 142896 218816
rect 142948 218804 142954 218816
rect 307110 218804 307116 218816
rect 142948 218776 307116 218804
rect 142948 218764 142954 218776
rect 307110 218764 307116 218776
rect 307168 218764 307174 218816
rect 50706 218696 50712 218748
rect 50764 218736 50770 218748
rect 311158 218736 311164 218748
rect 50764 218708 311164 218736
rect 50764 218696 50770 218708
rect 311158 218696 311164 218708
rect 311216 218696 311222 218748
rect 55030 217404 55036 217456
rect 55088 217444 55094 217456
rect 196710 217444 196716 217456
rect 55088 217416 196716 217444
rect 55088 217404 55094 217416
rect 196710 217404 196716 217416
rect 196768 217404 196774 217456
rect 67542 217336 67548 217388
rect 67600 217376 67606 217388
rect 251266 217376 251272 217388
rect 67600 217348 251272 217376
rect 67600 217336 67606 217348
rect 251266 217336 251272 217348
rect 251324 217336 251330 217388
rect 71038 217268 71044 217320
rect 71096 217308 71102 217320
rect 315390 217308 315396 217320
rect 71096 217280 315396 217308
rect 71096 217268 71102 217280
rect 315390 217268 315396 217280
rect 315448 217268 315454 217320
rect 304258 216696 304264 216708
rect 303908 216668 304264 216696
rect 122190 216588 122196 216640
rect 122248 216628 122254 216640
rect 303908 216628 303936 216668
rect 304258 216656 304264 216668
rect 304316 216696 304322 216708
rect 346670 216696 346676 216708
rect 304316 216668 346676 216696
rect 304316 216656 304322 216668
rect 346670 216656 346676 216668
rect 346728 216656 346734 216708
rect 122248 216600 303936 216628
rect 122248 216588 122254 216600
rect 93946 216520 93952 216572
rect 94004 216560 94010 216572
rect 146294 216560 146300 216572
rect 94004 216532 146300 216560
rect 94004 216520 94010 216532
rect 146294 216520 146300 216532
rect 146352 216520 146358 216572
rect 142982 216112 142988 216164
rect 143040 216152 143046 216164
rect 235258 216152 235264 216164
rect 143040 216124 235264 216152
rect 143040 216112 143046 216124
rect 235258 216112 235264 216124
rect 235316 216112 235322 216164
rect 50890 216044 50896 216096
rect 50948 216084 50954 216096
rect 162302 216084 162308 216096
rect 50948 216056 162308 216084
rect 50948 216044 50954 216056
rect 162302 216044 162308 216056
rect 162360 216044 162366 216096
rect 146294 215976 146300 216028
rect 146352 216016 146358 216028
rect 327074 216016 327080 216028
rect 146352 215988 327080 216016
rect 146352 215976 146358 215988
rect 327074 215976 327080 215988
rect 327132 215976 327138 216028
rect 74626 215908 74632 215960
rect 74684 215948 74690 215960
rect 280154 215948 280160 215960
rect 74684 215920 280160 215948
rect 74684 215908 74690 215920
rect 280154 215908 280160 215920
rect 280212 215908 280218 215960
rect 258074 215364 258080 215416
rect 258132 215404 258138 215416
rect 264238 215404 264244 215416
rect 258132 215376 264244 215404
rect 258132 215364 258138 215376
rect 264238 215364 264244 215376
rect 264296 215364 264302 215416
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 18598 215268 18604 215280
rect 3384 215240 18604 215268
rect 3384 215228 3390 215240
rect 18598 215228 18604 215240
rect 18656 215228 18662 215280
rect 103698 215228 103704 215280
rect 103756 215268 103762 215280
rect 164142 215268 164148 215280
rect 103756 215240 164148 215268
rect 103756 215228 103762 215240
rect 164142 215228 164148 215240
rect 164200 215228 164206 215280
rect 154022 214820 154028 214872
rect 154080 214860 154086 214872
rect 270586 214860 270592 214872
rect 154080 214832 270592 214860
rect 154080 214820 154086 214832
rect 270586 214820 270592 214832
rect 270644 214820 270650 214872
rect 50798 214752 50804 214804
rect 50856 214792 50862 214804
rect 211798 214792 211804 214804
rect 50856 214764 211804 214792
rect 50856 214752 50862 214764
rect 211798 214752 211804 214764
rect 211856 214752 211862 214804
rect 164142 214684 164148 214736
rect 164200 214724 164206 214736
rect 328454 214724 328460 214736
rect 164200 214696 328460 214724
rect 164200 214684 164206 214696
rect 328454 214684 328460 214696
rect 328512 214684 328518 214736
rect 57790 214616 57796 214668
rect 57848 214656 57854 214668
rect 250438 214656 250444 214668
rect 57848 214628 250444 214656
rect 57848 214616 57854 214628
rect 250438 214616 250444 214628
rect 250496 214616 250502 214668
rect 108942 214548 108948 214600
rect 109000 214588 109006 214600
rect 328638 214588 328644 214600
rect 109000 214560 328644 214588
rect 109000 214548 109006 214560
rect 328638 214548 328644 214560
rect 328696 214548 328702 214600
rect 84286 213868 84292 213920
rect 84344 213908 84350 213920
rect 133874 213908 133880 213920
rect 84344 213880 133880 213908
rect 84344 213868 84350 213880
rect 133874 213868 133880 213880
rect 133932 213908 133938 213920
rect 135162 213908 135168 213920
rect 133932 213880 135168 213908
rect 133932 213868 133938 213880
rect 135162 213868 135168 213880
rect 135220 213868 135226 213920
rect 147030 213324 147036 213376
rect 147088 213364 147094 213376
rect 259454 213364 259460 213376
rect 147088 213336 259460 213364
rect 147088 213324 147094 213336
rect 259454 213324 259460 213336
rect 259512 213324 259518 213376
rect 111794 213256 111800 213308
rect 111852 213296 111858 213308
rect 273346 213296 273352 213308
rect 111852 213268 273352 213296
rect 111852 213256 111858 213268
rect 273346 213256 273352 213268
rect 273404 213256 273410 213308
rect 25498 213188 25504 213240
rect 25556 213228 25562 213240
rect 83458 213228 83464 213240
rect 25556 213200 83464 213228
rect 25556 213188 25562 213200
rect 83458 213188 83464 213200
rect 83516 213188 83522 213240
rect 135162 213188 135168 213240
rect 135220 213228 135226 213240
rect 322934 213228 322940 213240
rect 135220 213200 322940 213228
rect 135220 213188 135226 213200
rect 322934 213188 322940 213200
rect 322992 213188 322998 213240
rect 137370 211964 137376 212016
rect 137428 212004 137434 212016
rect 224218 212004 224224 212016
rect 137428 211976 224224 212004
rect 137428 211964 137434 211976
rect 224218 211964 224224 211976
rect 224276 211964 224282 212016
rect 62022 211896 62028 211948
rect 62080 211936 62086 211948
rect 272058 211936 272064 211948
rect 62080 211908 272064 211936
rect 62080 211896 62086 211908
rect 272058 211896 272064 211908
rect 272116 211896 272122 211948
rect 78674 211828 78680 211880
rect 78732 211868 78738 211880
rect 328546 211868 328552 211880
rect 78732 211840 328552 211868
rect 78732 211828 78738 211840
rect 328546 211828 328552 211840
rect 328604 211828 328610 211880
rect 35710 211760 35716 211812
rect 35768 211800 35774 211812
rect 313918 211800 313924 211812
rect 35768 211772 313924 211800
rect 35768 211760 35774 211772
rect 313918 211760 313924 211772
rect 313976 211760 313982 211812
rect 289814 211148 289820 211200
rect 289872 211188 289878 211200
rect 296714 211188 296720 211200
rect 289872 211160 296720 211188
rect 289872 211148 289878 211160
rect 296714 211148 296720 211160
rect 296772 211148 296778 211200
rect 89714 210536 89720 210588
rect 89772 210576 89778 210588
rect 253934 210576 253940 210588
rect 89772 210548 253940 210576
rect 89772 210536 89778 210548
rect 253934 210536 253940 210548
rect 253992 210536 253998 210588
rect 129642 210468 129648 210520
rect 129700 210508 129706 210520
rect 335354 210508 335360 210520
rect 129700 210480 335360 210508
rect 129700 210468 129706 210480
rect 335354 210468 335360 210480
rect 335412 210468 335418 210520
rect 53466 210400 53472 210452
rect 53524 210440 53530 210452
rect 289078 210440 289084 210452
rect 53524 210412 289084 210440
rect 53524 210400 53530 210412
rect 289078 210400 289084 210412
rect 289136 210400 289142 210452
rect 43990 209720 43996 209772
rect 44048 209760 44054 209772
rect 327258 209760 327264 209772
rect 44048 209732 327264 209760
rect 44048 209720 44054 209732
rect 327258 209720 327264 209732
rect 327316 209720 327322 209772
rect 84194 209652 84200 209704
rect 84252 209692 84258 209704
rect 136634 209692 136640 209704
rect 84252 209664 136640 209692
rect 84252 209652 84258 209664
rect 136634 209652 136640 209664
rect 136692 209652 136698 209704
rect 126330 209176 126336 209228
rect 126388 209216 126394 209228
rect 233878 209216 233884 209228
rect 126388 209188 233884 209216
rect 126388 209176 126394 209188
rect 233878 209176 233884 209188
rect 233936 209176 233942 209228
rect 136634 209108 136640 209160
rect 136692 209148 136698 209160
rect 321646 209148 321652 209160
rect 136692 209120 321652 209148
rect 136692 209108 136698 209120
rect 321646 209108 321652 209120
rect 321704 209108 321710 209160
rect 86218 209040 86224 209092
rect 86276 209080 86282 209092
rect 277394 209080 277400 209092
rect 86276 209052 277400 209080
rect 86276 209040 86282 209052
rect 277394 209040 277400 209052
rect 277452 209040 277458 209092
rect 327258 209040 327264 209092
rect 327316 209080 327322 209092
rect 354674 209080 354680 209092
rect 327316 209052 354680 209080
rect 327316 209040 327322 209052
rect 354674 209040 354680 209052
rect 354732 209040 354738 209092
rect 114554 208292 114560 208344
rect 114612 208332 114618 208344
rect 169754 208332 169760 208344
rect 114612 208304 169760 208332
rect 114612 208292 114618 208304
rect 169754 208292 169760 208304
rect 169812 208292 169818 208344
rect 80054 208224 80060 208276
rect 80112 208264 80118 208276
rect 122834 208264 122840 208276
rect 80112 208236 122840 208264
rect 80112 208224 80118 208236
rect 122834 208224 122840 208236
rect 122892 208264 122898 208276
rect 124122 208264 124128 208276
rect 122892 208236 124128 208264
rect 122892 208224 122898 208236
rect 124122 208224 124128 208236
rect 124180 208224 124186 208276
rect 169754 207884 169760 207936
rect 169812 207924 169818 207936
rect 170858 207924 170864 207936
rect 169812 207896 170864 207924
rect 169812 207884 169818 207896
rect 170858 207884 170864 207896
rect 170916 207924 170922 207936
rect 186958 207924 186964 207936
rect 170916 207896 186964 207924
rect 170916 207884 170922 207896
rect 186958 207884 186964 207896
rect 187016 207884 187022 207936
rect 158070 207816 158076 207868
rect 158128 207856 158134 207868
rect 233970 207856 233976 207868
rect 158128 207828 233976 207856
rect 158128 207816 158134 207828
rect 233970 207816 233976 207828
rect 234028 207816 234034 207868
rect 245654 207816 245660 207868
rect 245712 207856 245718 207868
rect 308490 207856 308496 207868
rect 245712 207828 308496 207856
rect 245712 207816 245718 207828
rect 308490 207816 308496 207828
rect 308548 207816 308554 207868
rect 115934 207748 115940 207800
rect 115992 207788 115998 207800
rect 246298 207788 246304 207800
rect 115992 207760 246304 207788
rect 115992 207748 115998 207760
rect 246298 207748 246304 207760
rect 246356 207748 246362 207800
rect 124122 207680 124128 207732
rect 124180 207720 124186 207732
rect 330110 207720 330116 207732
rect 124180 207692 330116 207720
rect 124180 207680 124186 207692
rect 330110 207680 330116 207692
rect 330168 207680 330174 207732
rect 54938 207612 54944 207664
rect 54996 207652 55002 207664
rect 318150 207652 318156 207664
rect 54996 207624 318156 207652
rect 54996 207612 55002 207624
rect 318150 207612 318156 207624
rect 318208 207612 318214 207664
rect 574738 206932 574744 206984
rect 574796 206972 574802 206984
rect 579890 206972 579896 206984
rect 574796 206944 579896 206972
rect 574796 206932 574802 206944
rect 579890 206932 579896 206944
rect 579948 206932 579954 206984
rect 248414 206592 248420 206644
rect 248472 206632 248478 206644
rect 287698 206632 287704 206644
rect 248472 206604 287704 206632
rect 248472 206592 248478 206604
rect 287698 206592 287704 206604
rect 287756 206592 287762 206644
rect 149974 206524 149980 206576
rect 150032 206564 150038 206576
rect 270678 206564 270684 206576
rect 150032 206536 270684 206564
rect 150032 206524 150038 206536
rect 270678 206524 270684 206536
rect 270736 206524 270742 206576
rect 168006 206456 168012 206508
rect 168064 206496 168070 206508
rect 345014 206496 345020 206508
rect 168064 206468 345020 206496
rect 168064 206456 168070 206468
rect 345014 206456 345020 206468
rect 345072 206456 345078 206508
rect 66162 206388 66168 206440
rect 66220 206428 66226 206440
rect 251358 206428 251364 206440
rect 66220 206400 251364 206428
rect 66220 206388 66226 206400
rect 251358 206388 251364 206400
rect 251416 206388 251422 206440
rect 274634 206388 274640 206440
rect 274692 206428 274698 206440
rect 293218 206428 293224 206440
rect 274692 206400 293224 206428
rect 274692 206388 274698 206400
rect 293218 206388 293224 206400
rect 293276 206388 293282 206440
rect 133138 206320 133144 206372
rect 133196 206360 133202 206372
rect 350626 206360 350632 206372
rect 133196 206332 350632 206360
rect 133196 206320 133202 206332
rect 350626 206320 350632 206332
rect 350684 206320 350690 206372
rect 104250 206252 104256 206304
rect 104308 206292 104314 206304
rect 339586 206292 339592 206304
rect 104308 206264 339592 206292
rect 104308 206252 104314 206264
rect 339586 206252 339592 206264
rect 339644 206252 339650 206304
rect 96430 205572 96436 205624
rect 96488 205612 96494 205624
rect 146202 205612 146208 205624
rect 96488 205584 146208 205612
rect 96488 205572 96494 205584
rect 146202 205572 146208 205584
rect 146260 205572 146266 205624
rect 146202 205028 146208 205080
rect 146260 205068 146266 205080
rect 346486 205068 346492 205080
rect 146260 205040 346492 205068
rect 146260 205028 146266 205040
rect 346486 205028 346492 205040
rect 346544 205028 346550 205080
rect 48038 204960 48044 205012
rect 48096 205000 48102 205012
rect 278958 205000 278964 205012
rect 48096 204972 278964 205000
rect 48096 204960 48102 204972
rect 278958 204960 278964 204972
rect 279016 204960 279022 205012
rect 74534 204892 74540 204944
rect 74592 204932 74598 204944
rect 343726 204932 343732 204944
rect 74592 204904 343732 204932
rect 74592 204892 74598 204904
rect 343726 204892 343732 204904
rect 343784 204892 343790 204944
rect 146938 203804 146944 203856
rect 146996 203844 147002 203856
rect 264974 203844 264980 203856
rect 146996 203816 264980 203844
rect 146996 203804 147002 203816
rect 264974 203804 264980 203816
rect 265032 203804 265038 203856
rect 133230 203736 133236 203788
rect 133288 203776 133294 203788
rect 267826 203776 267832 203788
rect 133288 203748 267832 203776
rect 133288 203736 133294 203748
rect 267826 203736 267832 203748
rect 267884 203736 267890 203788
rect 110414 203668 110420 203720
rect 110472 203708 110478 203720
rect 249794 203708 249800 203720
rect 110472 203680 249800 203708
rect 110472 203668 110478 203680
rect 249794 203668 249800 203680
rect 249852 203668 249858 203720
rect 271874 203668 271880 203720
rect 271932 203708 271938 203720
rect 294046 203708 294052 203720
rect 271932 203680 294052 203708
rect 271932 203668 271938 203680
rect 294046 203668 294052 203680
rect 294104 203668 294110 203720
rect 92474 203600 92480 203652
rect 92532 203640 92538 203652
rect 242158 203640 242164 203652
rect 92532 203612 242164 203640
rect 92532 203600 92538 203612
rect 242158 203600 242164 203612
rect 242216 203600 242222 203652
rect 281534 203600 281540 203652
rect 281592 203640 281598 203652
rect 342346 203640 342352 203652
rect 281592 203612 342352 203640
rect 281592 203600 281598 203612
rect 342346 203600 342352 203612
rect 342404 203600 342410 203652
rect 72418 203532 72424 203584
rect 72476 203572 72482 203584
rect 325878 203572 325884 203584
rect 72476 203544 325884 203572
rect 72476 203532 72482 203544
rect 325878 203532 325884 203544
rect 325936 203532 325942 203584
rect 119982 202240 119988 202292
rect 120040 202280 120046 202292
rect 329834 202280 329840 202292
rect 120040 202252 329840 202280
rect 120040 202240 120046 202252
rect 329834 202240 329840 202252
rect 329892 202240 329898 202292
rect 66070 202172 66076 202224
rect 66128 202212 66134 202224
rect 278866 202212 278872 202224
rect 66128 202184 278872 202212
rect 66128 202172 66134 202184
rect 278866 202172 278872 202184
rect 278924 202172 278930 202224
rect 99374 202104 99380 202156
rect 99432 202144 99438 202156
rect 327350 202144 327356 202156
rect 99432 202116 327356 202144
rect 99432 202104 99438 202116
rect 327350 202104 327356 202116
rect 327408 202104 327414 202156
rect 158162 200880 158168 200932
rect 158220 200920 158226 200932
rect 256970 200920 256976 200932
rect 158220 200892 256976 200920
rect 158220 200880 158226 200892
rect 256970 200880 256976 200892
rect 257028 200880 257034 200932
rect 131850 200812 131856 200864
rect 131908 200852 131914 200864
rect 318242 200852 318248 200864
rect 131908 200824 318248 200852
rect 131908 200812 131914 200824
rect 318242 200812 318248 200824
rect 318300 200812 318306 200864
rect 153930 200744 153936 200796
rect 153988 200784 153994 200796
rect 351914 200784 351920 200796
rect 153988 200756 351920 200784
rect 153988 200744 153994 200756
rect 351914 200744 351920 200756
rect 351972 200744 351978 200796
rect 157978 199588 157984 199640
rect 158036 199628 158042 199640
rect 246390 199628 246396 199640
rect 158036 199600 246396 199628
rect 158036 199588 158042 199600
rect 246390 199588 246396 199600
rect 246448 199588 246454 199640
rect 134518 199520 134524 199572
rect 134576 199560 134582 199572
rect 242250 199560 242256 199572
rect 134576 199532 242256 199560
rect 134576 199520 134582 199532
rect 242250 199520 242256 199532
rect 242308 199520 242314 199572
rect 69290 199452 69296 199504
rect 69348 199492 69354 199504
rect 248506 199492 248512 199504
rect 69348 199464 248512 199492
rect 69348 199452 69354 199464
rect 248506 199452 248512 199464
rect 248564 199452 248570 199504
rect 93762 199384 93768 199436
rect 93820 199424 93826 199436
rect 347866 199424 347872 199436
rect 93820 199396 347872 199424
rect 93820 199384 93826 199396
rect 347866 199384 347872 199396
rect 347924 199384 347930 199436
rect 160830 198160 160836 198212
rect 160888 198200 160894 198212
rect 266354 198200 266360 198212
rect 160888 198172 266360 198200
rect 160888 198160 160894 198172
rect 266354 198160 266360 198172
rect 266412 198160 266418 198212
rect 138658 198092 138664 198144
rect 138716 198132 138722 198144
rect 276106 198132 276112 198144
rect 138716 198104 276112 198132
rect 138716 198092 138722 198104
rect 276106 198092 276112 198104
rect 276164 198092 276170 198144
rect 126238 198024 126244 198076
rect 126296 198064 126302 198076
rect 311250 198064 311256 198076
rect 126296 198036 311256 198064
rect 126296 198024 126302 198036
rect 311250 198024 311256 198036
rect 311308 198024 311314 198076
rect 77938 197956 77944 198008
rect 77996 197996 78002 198008
rect 330018 197996 330024 198008
rect 77996 197968 330024 197996
rect 77996 197956 78002 197968
rect 330018 197956 330024 197968
rect 330076 197956 330082 198008
rect 144362 196868 144368 196920
rect 144420 196908 144426 196920
rect 262398 196908 262404 196920
rect 144420 196880 262404 196908
rect 144420 196868 144426 196880
rect 262398 196868 262404 196880
rect 262456 196868 262462 196920
rect 222838 196800 222844 196852
rect 222896 196840 222902 196852
rect 354766 196840 354772 196852
rect 222896 196812 354772 196840
rect 222896 196800 222902 196812
rect 354766 196800 354772 196812
rect 354824 196800 354830 196852
rect 96614 196732 96620 196784
rect 96672 196772 96678 196784
rect 249058 196772 249064 196784
rect 96672 196744 249064 196772
rect 96672 196732 96678 196744
rect 249058 196732 249064 196744
rect 249116 196732 249122 196784
rect 63126 196664 63132 196716
rect 63184 196704 63190 196716
rect 271966 196704 271972 196716
rect 63184 196676 271972 196704
rect 63184 196664 63190 196676
rect 271966 196664 271972 196676
rect 272024 196664 272030 196716
rect 56410 196596 56416 196648
rect 56468 196636 56474 196648
rect 276014 196636 276020 196648
rect 56468 196608 276020 196636
rect 56468 196596 56474 196608
rect 276014 196596 276020 196608
rect 276072 196596 276078 196648
rect 138842 195440 138848 195492
rect 138900 195480 138906 195492
rect 239490 195480 239496 195492
rect 138900 195452 239496 195480
rect 138900 195440 138906 195452
rect 239490 195440 239496 195452
rect 239548 195440 239554 195492
rect 91738 195372 91744 195424
rect 91796 195412 91802 195424
rect 246482 195412 246488 195424
rect 91796 195384 246488 195412
rect 91796 195372 91802 195384
rect 246482 195372 246488 195384
rect 246540 195372 246546 195424
rect 163498 195304 163504 195356
rect 163556 195344 163562 195356
rect 334250 195344 334256 195356
rect 163556 195316 334256 195344
rect 163556 195304 163562 195316
rect 334250 195304 334256 195316
rect 334308 195304 334314 195356
rect 160738 195236 160744 195288
rect 160796 195276 160802 195288
rect 582466 195276 582472 195288
rect 160796 195248 582472 195276
rect 160796 195236 160802 195248
rect 582466 195236 582472 195248
rect 582524 195236 582530 195288
rect 99282 194012 99288 194064
rect 99340 194052 99346 194064
rect 162394 194052 162400 194064
rect 99340 194024 162400 194052
rect 99340 194012 99346 194024
rect 162394 194012 162400 194024
rect 162452 194012 162458 194064
rect 124950 193944 124956 193996
rect 125008 193984 125014 193996
rect 231118 193984 231124 193996
rect 125008 193956 231124 193984
rect 125008 193944 125014 193956
rect 231118 193944 231124 193956
rect 231176 193944 231182 193996
rect 144270 193876 144276 193928
rect 144328 193916 144334 193928
rect 266446 193916 266452 193928
rect 144328 193888 266452 193916
rect 144328 193876 144334 193888
rect 266446 193876 266452 193888
rect 266504 193876 266510 193928
rect 140130 193808 140136 193860
rect 140188 193848 140194 193860
rect 340966 193848 340972 193860
rect 140188 193820 340972 193848
rect 140188 193808 140194 193820
rect 340966 193808 340972 193820
rect 341024 193808 341030 193860
rect 227714 192720 227720 192772
rect 227772 192760 227778 192772
rect 346394 192760 346400 192772
rect 227772 192732 346400 192760
rect 227772 192720 227778 192732
rect 346394 192720 346400 192732
rect 346452 192720 346458 192772
rect 100754 192652 100760 192704
rect 100812 192692 100818 192704
rect 254026 192692 254032 192704
rect 100812 192664 254032 192692
rect 100812 192652 100818 192664
rect 254026 192652 254032 192664
rect 254084 192652 254090 192704
rect 77294 192584 77300 192636
rect 77352 192624 77358 192636
rect 252646 192624 252652 192636
rect 77352 192596 252652 192624
rect 77352 192584 77358 192596
rect 252646 192584 252652 192596
rect 252704 192584 252710 192636
rect 104158 192516 104164 192568
rect 104216 192556 104222 192568
rect 321554 192556 321560 192568
rect 104216 192528 321560 192556
rect 104216 192516 104222 192528
rect 321554 192516 321560 192528
rect 321612 192516 321618 192568
rect 49602 192448 49608 192500
rect 49660 192488 49666 192500
rect 269206 192488 269212 192500
rect 49660 192460 269212 192488
rect 49660 192448 49666 192460
rect 269206 192448 269212 192460
rect 269264 192448 269270 192500
rect 124858 191360 124864 191412
rect 124916 191400 124922 191412
rect 185578 191400 185584 191412
rect 124916 191372 185584 191400
rect 124916 191360 124922 191372
rect 185578 191360 185584 191372
rect 185636 191360 185642 191412
rect 204162 191360 204168 191412
rect 204220 191400 204226 191412
rect 220814 191400 220820 191412
rect 204220 191372 220820 191400
rect 204220 191360 204226 191372
rect 220814 191360 220820 191372
rect 220872 191360 220878 191412
rect 136082 191292 136088 191344
rect 136140 191332 136146 191344
rect 242342 191332 242348 191344
rect 136140 191304 242348 191332
rect 136140 191292 136146 191304
rect 242342 191292 242348 191304
rect 242400 191292 242406 191344
rect 148502 191224 148508 191276
rect 148560 191264 148566 191276
rect 255406 191264 255412 191276
rect 148560 191236 255412 191264
rect 148560 191224 148566 191236
rect 255406 191224 255412 191236
rect 255464 191224 255470 191276
rect 53742 191156 53748 191208
rect 53800 191196 53806 191208
rect 259546 191196 259552 191208
rect 53800 191168 259552 191196
rect 53800 191156 53806 191168
rect 259546 191156 259552 191168
rect 259604 191156 259610 191208
rect 264330 191156 264336 191208
rect 264388 191196 264394 191208
rect 342530 191196 342536 191208
rect 264388 191168 342536 191196
rect 264388 191156 264394 191168
rect 342530 191156 342536 191168
rect 342588 191156 342594 191208
rect 70394 191088 70400 191140
rect 70452 191128 70458 191140
rect 315482 191128 315488 191140
rect 70452 191100 315488 191128
rect 70452 191088 70458 191100
rect 315482 191088 315488 191100
rect 315540 191088 315546 191140
rect 214558 190068 214564 190120
rect 214616 190108 214622 190120
rect 274818 190108 274824 190120
rect 214616 190080 274824 190108
rect 214616 190068 214622 190080
rect 274818 190068 274824 190080
rect 274876 190068 274882 190120
rect 160002 190000 160008 190052
rect 160060 190040 160066 190052
rect 196618 190040 196624 190052
rect 160060 190012 196624 190040
rect 160060 190000 160066 190012
rect 196618 190000 196624 190012
rect 196676 190000 196682 190052
rect 237374 190000 237380 190052
rect 237432 190040 237438 190052
rect 340874 190040 340880 190052
rect 237432 190012 340880 190040
rect 237432 190000 237438 190012
rect 340874 190000 340880 190012
rect 340932 190000 340938 190052
rect 153838 189932 153844 189984
rect 153896 189972 153902 189984
rect 258166 189972 258172 189984
rect 153896 189944 258172 189972
rect 153896 189932 153902 189944
rect 258166 189932 258172 189944
rect 258224 189932 258230 189984
rect 102134 189864 102140 189916
rect 102192 189904 102198 189916
rect 249978 189904 249984 189916
rect 102192 189876 249984 189904
rect 102192 189864 102198 189876
rect 249978 189864 249984 189876
rect 250036 189864 250042 189916
rect 18598 189796 18604 189848
rect 18656 189836 18662 189848
rect 109034 189836 109040 189848
rect 18656 189808 109040 189836
rect 18656 189796 18662 189808
rect 109034 189796 109040 189808
rect 109092 189796 109098 189848
rect 169386 189796 169392 189848
rect 169444 189836 169450 189848
rect 341058 189836 341064 189848
rect 169444 189808 341064 189836
rect 169444 189796 169450 189808
rect 341058 189796 341064 189808
rect 341116 189796 341122 189848
rect 88242 189728 88248 189780
rect 88300 189768 88306 189780
rect 327258 189768 327264 189780
rect 88300 189740 327264 189768
rect 88300 189728 88306 189740
rect 327258 189728 327264 189740
rect 327316 189728 327322 189780
rect 106182 189116 106188 189168
rect 106240 189156 106246 189168
rect 169202 189156 169208 189168
rect 106240 189128 169208 189156
rect 106240 189116 106246 189128
rect 169202 189116 169208 189128
rect 169260 189116 169266 189168
rect 134518 189048 134524 189100
rect 134576 189088 134582 189100
rect 214650 189088 214656 189100
rect 134576 189060 214656 189088
rect 134576 189048 134582 189060
rect 214650 189048 214656 189060
rect 214708 189048 214714 189100
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 59998 189020 60004 189032
rect 3476 188992 60004 189020
rect 3476 188980 3482 188992
rect 59998 188980 60004 188992
rect 60056 188980 60062 189032
rect 140038 188436 140044 188488
rect 140096 188476 140102 188488
rect 263686 188476 263692 188488
rect 140096 188448 263692 188476
rect 140096 188436 140102 188448
rect 263686 188436 263692 188448
rect 263744 188436 263750 188488
rect 127618 188368 127624 188420
rect 127676 188408 127682 188420
rect 269298 188408 269304 188420
rect 127676 188380 269304 188408
rect 127676 188368 127682 188380
rect 269298 188368 269304 188380
rect 269356 188368 269362 188420
rect 66990 188300 66996 188352
rect 67048 188340 67054 188352
rect 319530 188340 319536 188352
rect 67048 188312 319536 188340
rect 67048 188300 67054 188312
rect 319530 188300 319536 188312
rect 319588 188300 319594 188352
rect 102042 187688 102048 187740
rect 102100 187728 102106 187740
rect 184198 187728 184204 187740
rect 102100 187700 184204 187728
rect 102100 187688 102106 187700
rect 184198 187688 184204 187700
rect 184256 187688 184262 187740
rect 157150 187212 157156 187264
rect 157208 187252 157214 187264
rect 198090 187252 198096 187264
rect 157208 187224 198096 187252
rect 157208 187212 157214 187224
rect 198090 187212 198096 187224
rect 198148 187212 198154 187264
rect 131758 187144 131764 187196
rect 131816 187184 131822 187196
rect 267734 187184 267740 187196
rect 131816 187156 267740 187184
rect 131816 187144 131822 187156
rect 267734 187144 267740 187156
rect 267792 187144 267798 187196
rect 173158 187076 173164 187128
rect 173216 187116 173222 187128
rect 324498 187116 324504 187128
rect 173216 187088 324504 187116
rect 173216 187076 173222 187088
rect 324498 187076 324504 187088
rect 324556 187076 324562 187128
rect 49510 187008 49516 187060
rect 49568 187048 49574 187060
rect 256786 187048 256792 187060
rect 49568 187020 256792 187048
rect 49568 187008 49574 187020
rect 256786 187008 256792 187020
rect 256844 187008 256850 187060
rect 96522 186940 96528 186992
rect 96580 186980 96586 186992
rect 321830 186980 321836 186992
rect 96580 186952 321836 186980
rect 96580 186940 96586 186952
rect 321830 186940 321836 186952
rect 321888 186940 321894 186992
rect 323670 186940 323676 186992
rect 323728 186980 323734 186992
rect 332686 186980 332692 186992
rect 323728 186952 332692 186980
rect 323728 186940 323734 186952
rect 332686 186940 332692 186952
rect 332744 186940 332750 186992
rect 132402 186396 132408 186448
rect 132460 186436 132466 186448
rect 167914 186436 167920 186448
rect 132460 186408 167920 186436
rect 132460 186396 132466 186408
rect 167914 186396 167920 186408
rect 167972 186396 167978 186448
rect 104802 186328 104808 186380
rect 104860 186368 104866 186380
rect 173250 186368 173256 186380
rect 104860 186340 173256 186368
rect 104860 186328 104866 186340
rect 173250 186328 173256 186340
rect 173308 186328 173314 186380
rect 196710 185784 196716 185836
rect 196768 185824 196774 185836
rect 259638 185824 259644 185836
rect 196768 185796 259644 185824
rect 196768 185784 196774 185796
rect 259638 185784 259644 185796
rect 259696 185784 259702 185836
rect 141418 185716 141424 185768
rect 141476 185756 141482 185768
rect 255590 185756 255596 185768
rect 141476 185728 255596 185756
rect 141476 185716 141482 185728
rect 255590 185716 255596 185728
rect 255648 185716 255654 185768
rect 148410 185648 148416 185700
rect 148468 185688 148474 185700
rect 318426 185688 318432 185700
rect 148468 185660 318432 185688
rect 148468 185648 148474 185660
rect 318426 185648 318432 185660
rect 318484 185648 318490 185700
rect 73798 185580 73804 185632
rect 73856 185620 73862 185632
rect 321278 185620 321284 185632
rect 73856 185592 321284 185620
rect 73856 185580 73862 185592
rect 321278 185580 321284 185592
rect 321336 185580 321342 185632
rect 100662 184968 100668 185020
rect 100720 185008 100726 185020
rect 170398 185008 170404 185020
rect 100720 184980 170404 185008
rect 100720 184968 100726 184980
rect 170398 184968 170404 184980
rect 170456 184968 170462 185020
rect 125502 184900 125508 184952
rect 125560 184940 125566 184952
rect 214926 184940 214932 184952
rect 125560 184912 214932 184940
rect 125560 184900 125566 184912
rect 214926 184900 214932 184912
rect 214984 184900 214990 184952
rect 155862 184492 155868 184544
rect 155920 184532 155926 184544
rect 192570 184532 192576 184544
rect 155920 184504 192576 184532
rect 155920 184492 155926 184504
rect 192570 184492 192576 184504
rect 192628 184492 192634 184544
rect 203518 184492 203524 184544
rect 203576 184532 203582 184544
rect 259730 184532 259736 184544
rect 203576 184504 259736 184532
rect 203576 184492 203582 184504
rect 259730 184492 259736 184504
rect 259788 184492 259794 184544
rect 149790 184424 149796 184476
rect 149848 184464 149854 184476
rect 274726 184464 274732 184476
rect 149848 184436 274732 184464
rect 149848 184424 149854 184436
rect 274726 184424 274732 184436
rect 274784 184424 274790 184476
rect 64690 184356 64696 184408
rect 64748 184396 64754 184408
rect 254210 184396 254216 184408
rect 64748 184368 254216 184396
rect 64748 184356 64754 184368
rect 254210 184356 254216 184368
rect 254268 184356 254274 184408
rect 319438 184356 319444 184408
rect 319496 184396 319502 184408
rect 332778 184396 332784 184408
rect 319496 184368 332784 184396
rect 319496 184356 319502 184368
rect 332778 184356 332784 184368
rect 332836 184356 332842 184408
rect 111150 184288 111156 184340
rect 111208 184328 111214 184340
rect 339770 184328 339776 184340
rect 111208 184300 339776 184328
rect 111208 184288 111214 184300
rect 339770 184288 339776 184300
rect 339828 184288 339834 184340
rect 69658 184220 69664 184272
rect 69716 184260 69722 184272
rect 338390 184260 338396 184272
rect 69716 184232 338396 184260
rect 69716 184220 69722 184232
rect 338390 184220 338396 184232
rect 338448 184220 338454 184272
rect 75178 184152 75184 184204
rect 75236 184192 75242 184204
rect 347958 184192 347964 184204
rect 75236 184164 347964 184192
rect 75236 184152 75242 184164
rect 347958 184152 347964 184164
rect 348016 184152 348022 184204
rect 157242 182996 157248 183048
rect 157300 183036 157306 183048
rect 191098 183036 191104 183048
rect 157300 183008 191104 183036
rect 157300 182996 157306 183008
rect 191098 182996 191104 183008
rect 191156 182996 191162 183048
rect 224218 182996 224224 183048
rect 224276 183036 224282 183048
rect 260926 183036 260932 183048
rect 224276 183008 260932 183036
rect 224276 182996 224282 183008
rect 260926 182996 260932 183008
rect 260984 182996 260990 183048
rect 162210 182928 162216 182980
rect 162268 182968 162274 182980
rect 338206 182968 338212 182980
rect 162268 182940 338212 182968
rect 162268 182928 162274 182940
rect 338206 182928 338212 182940
rect 338264 182928 338270 182980
rect 122098 182860 122104 182912
rect 122156 182900 122162 182912
rect 345198 182900 345204 182912
rect 122156 182872 345204 182900
rect 122156 182860 122162 182872
rect 345198 182860 345204 182872
rect 345256 182860 345262 182912
rect 73062 182792 73068 182844
rect 73120 182832 73126 182844
rect 336826 182832 336832 182844
rect 73120 182804 336832 182832
rect 73120 182792 73126 182804
rect 336826 182792 336832 182804
rect 336884 182792 336890 182844
rect 118418 182180 118424 182232
rect 118476 182220 118482 182232
rect 167822 182220 167828 182232
rect 118476 182192 167828 182220
rect 118476 182180 118482 182192
rect 167822 182180 167828 182192
rect 167880 182180 167886 182232
rect 240778 181704 240784 181756
rect 240836 181744 240842 181756
rect 262214 181744 262220 181756
rect 240836 181716 262220 181744
rect 240836 181704 240842 181716
rect 262214 181704 262220 181716
rect 262272 181704 262278 181756
rect 232498 181636 232504 181688
rect 232556 181676 232562 181688
rect 258258 181676 258264 181688
rect 232556 181648 258264 181676
rect 232556 181636 232562 181648
rect 258258 181636 258264 181648
rect 258316 181636 258322 181688
rect 318058 181636 318064 181688
rect 318116 181676 318122 181688
rect 338298 181676 338304 181688
rect 318116 181648 338304 181676
rect 318116 181636 318122 181648
rect 338298 181636 338304 181648
rect 338356 181636 338362 181688
rect 94038 181568 94044 181620
rect 94096 181608 94102 181620
rect 249886 181608 249892 181620
rect 94096 181580 249892 181608
rect 94096 181568 94102 181580
rect 249886 181568 249892 181580
rect 249944 181568 249950 181620
rect 289078 181568 289084 181620
rect 289136 181608 289142 181620
rect 334066 181608 334072 181620
rect 289136 181580 334072 181608
rect 289136 181568 289142 181580
rect 334066 181568 334072 181580
rect 334124 181568 334130 181620
rect 167730 181500 167736 181552
rect 167788 181540 167794 181552
rect 345106 181540 345112 181552
rect 167788 181512 345112 181540
rect 167788 181500 167794 181512
rect 345106 181500 345112 181512
rect 345164 181500 345170 181552
rect 41230 181432 41236 181484
rect 41288 181472 41294 181484
rect 313826 181472 313832 181484
rect 41288 181444 313832 181472
rect 41288 181432 41294 181444
rect 313826 181432 313832 181444
rect 313884 181432 313890 181484
rect 314562 181432 314568 181484
rect 314620 181472 314626 181484
rect 336734 181472 336740 181484
rect 314620 181444 336740 181472
rect 314620 181432 314626 181444
rect 336734 181432 336740 181444
rect 336792 181432 336798 181484
rect 133598 180888 133604 180940
rect 133656 180928 133662 180940
rect 164326 180928 164332 180940
rect 133656 180900 164332 180928
rect 133656 180888 133662 180900
rect 164326 180888 164332 180900
rect 164384 180888 164390 180940
rect 122006 180820 122012 180872
rect 122064 180860 122070 180872
rect 211982 180860 211988 180872
rect 122064 180832 211988 180860
rect 122064 180820 122070 180832
rect 211982 180820 211988 180832
rect 212040 180820 212046 180872
rect 244918 180344 244924 180396
rect 244976 180384 244982 180396
rect 255498 180384 255504 180396
rect 244976 180356 255504 180384
rect 244976 180344 244982 180356
rect 255498 180344 255504 180356
rect 255556 180344 255562 180396
rect 242158 180276 242164 180328
rect 242216 180316 242222 180328
rect 256878 180316 256884 180328
rect 242216 180288 256884 180316
rect 242216 180276 242222 180288
rect 256878 180276 256884 180288
rect 256936 180276 256942 180328
rect 244274 180208 244280 180260
rect 244332 180248 244338 180260
rect 270494 180248 270500 180260
rect 244332 180220 270500 180248
rect 244332 180208 244338 180220
rect 270494 180208 270500 180220
rect 270552 180208 270558 180260
rect 167638 180140 167644 180192
rect 167696 180180 167702 180192
rect 196710 180180 196716 180192
rect 167696 180152 196716 180180
rect 167696 180140 167702 180152
rect 196710 180140 196716 180152
rect 196768 180140 196774 180192
rect 233970 180140 233976 180192
rect 234028 180180 234034 180192
rect 260834 180180 260840 180192
rect 234028 180152 260840 180180
rect 234028 180140 234034 180152
rect 260834 180140 260840 180152
rect 260892 180140 260898 180192
rect 64782 180072 64788 180124
rect 64840 180112 64846 180124
rect 251450 180112 251456 180124
rect 64840 180084 251456 180112
rect 64840 180072 64846 180084
rect 251450 180072 251456 180084
rect 251508 180072 251514 180124
rect 315298 180072 315304 180124
rect 315356 180112 315362 180124
rect 341150 180112 341156 180124
rect 315356 180084 341156 180112
rect 315356 180072 315362 180084
rect 341150 180072 341156 180084
rect 341208 180072 341214 180124
rect 123018 179596 123024 179648
rect 123076 179636 123082 179648
rect 166350 179636 166356 179648
rect 123076 179608 166356 179636
rect 123076 179596 123082 179608
rect 166350 179596 166356 179608
rect 166408 179596 166414 179648
rect 120994 179528 121000 179580
rect 121052 179568 121058 179580
rect 167730 179568 167736 179580
rect 121052 179540 167736 179568
rect 121052 179528 121058 179540
rect 167730 179528 167736 179540
rect 167788 179528 167794 179580
rect 128170 179460 128176 179512
rect 128228 179500 128234 179512
rect 214098 179500 214104 179512
rect 128228 179472 214104 179500
rect 128228 179460 128234 179472
rect 214098 179460 214104 179472
rect 214156 179460 214162 179512
rect 114278 179392 114284 179444
rect 114336 179432 114342 179444
rect 209038 179432 209044 179444
rect 114336 179404 209044 179432
rect 114336 179392 114342 179404
rect 209038 179392 209044 179404
rect 209096 179392 209102 179444
rect 172146 179324 172152 179376
rect 172204 179364 172210 179376
rect 346302 179364 346308 179376
rect 172204 179336 346308 179364
rect 172204 179324 172210 179336
rect 346302 179324 346308 179336
rect 346360 179324 346366 179376
rect 169018 179256 169024 179308
rect 169076 179296 169082 179308
rect 342622 179296 342628 179308
rect 169076 179268 342628 179296
rect 169076 179256 169082 179268
rect 342622 179256 342628 179268
rect 342680 179256 342686 179308
rect 242342 178780 242348 178832
rect 242400 178820 242406 178832
rect 258442 178820 258448 178832
rect 242400 178792 258448 178820
rect 242400 178780 242406 178792
rect 258442 178780 258448 178792
rect 258500 178780 258506 178832
rect 211798 178712 211804 178764
rect 211856 178752 211862 178764
rect 258074 178752 258080 178764
rect 211856 178724 258080 178752
rect 211856 178712 211862 178724
rect 258074 178712 258080 178724
rect 258132 178712 258138 178764
rect 311250 178712 311256 178764
rect 311308 178752 311314 178764
rect 332686 178752 332692 178764
rect 311308 178724 332692 178752
rect 311308 178712 311314 178724
rect 332686 178712 332692 178724
rect 332744 178712 332750 178764
rect 138750 178644 138756 178696
rect 138808 178684 138814 178696
rect 252554 178684 252560 178696
rect 138808 178656 252560 178684
rect 138808 178644 138814 178656
rect 252554 178644 252560 178656
rect 252612 178644 252618 178696
rect 312538 178644 312544 178696
rect 312596 178684 312602 178696
rect 338114 178684 338120 178696
rect 312596 178656 338120 178684
rect 312596 178644 312602 178656
rect 338114 178644 338120 178656
rect 338172 178644 338178 178696
rect 112438 178236 112444 178288
rect 112496 178276 112502 178288
rect 211890 178276 211896 178288
rect 112496 178248 211896 178276
rect 112496 178236 112502 178248
rect 211890 178236 211896 178248
rect 211948 178236 211954 178288
rect 130746 178168 130752 178220
rect 130804 178208 130810 178220
rect 165522 178208 165528 178220
rect 130804 178180 165528 178208
rect 130804 178168 130810 178180
rect 165522 178168 165528 178180
rect 165580 178168 165586 178220
rect 148226 178100 148232 178152
rect 148284 178140 148290 178152
rect 214558 178140 214564 178152
rect 148284 178112 214564 178140
rect 148284 178100 148290 178112
rect 214558 178100 214564 178112
rect 214616 178100 214622 178152
rect 159910 178032 159916 178084
rect 159968 178072 159974 178084
rect 167638 178072 167644 178084
rect 159968 178044 167644 178072
rect 159968 178032 159974 178044
rect 167638 178032 167644 178044
rect 167696 178032 167702 178084
rect 289078 178032 289084 178084
rect 289136 178072 289142 178084
rect 316034 178072 316040 178084
rect 289136 178044 316040 178072
rect 289136 178032 289142 178044
rect 316034 178032 316040 178044
rect 316092 178032 316098 178084
rect 52546 177964 52552 178016
rect 52604 178004 52610 178016
rect 120074 178004 120080 178016
rect 52604 177976 120080 178004
rect 52604 177964 52610 177976
rect 120074 177964 120080 177976
rect 120132 177964 120138 178016
rect 242250 177964 242256 178016
rect 242308 178004 242314 178016
rect 249334 178004 249340 178016
rect 242308 177976 249340 178004
rect 242308 177964 242314 177976
rect 249334 177964 249340 177976
rect 249392 177964 249398 178016
rect 109954 177896 109960 177948
rect 110012 177936 110018 177948
rect 134518 177936 134524 177948
rect 110012 177908 134524 177936
rect 110012 177896 110018 177908
rect 134518 177896 134524 177908
rect 134576 177896 134582 177948
rect 239490 177556 239496 177608
rect 239548 177596 239554 177608
rect 256694 177596 256700 177608
rect 239548 177568 256700 177596
rect 239548 177556 239554 177568
rect 256694 177556 256700 177568
rect 256752 177556 256758 177608
rect 246482 177488 246488 177540
rect 246540 177528 246546 177540
rect 267918 177528 267924 177540
rect 246540 177500 267924 177528
rect 246540 177488 246546 177500
rect 267918 177488 267924 177500
rect 267976 177488 267982 177540
rect 315482 177488 315488 177540
rect 315540 177528 315546 177540
rect 331398 177528 331404 177540
rect 315540 177500 331404 177528
rect 315540 177488 315546 177500
rect 331398 177488 331404 177500
rect 331456 177488 331462 177540
rect 233878 177420 233884 177472
rect 233936 177460 233942 177472
rect 258350 177460 258356 177472
rect 233936 177432 258356 177460
rect 233936 177420 233942 177432
rect 258350 177420 258356 177432
rect 258408 177420 258414 177472
rect 311158 177420 311164 177472
rect 311216 177460 311222 177472
rect 331214 177460 331220 177472
rect 311216 177432 331220 177460
rect 311216 177420 311222 177432
rect 331214 177420 331220 177432
rect 331272 177420 331278 177472
rect 220078 177352 220084 177404
rect 220136 177392 220142 177404
rect 262306 177392 262312 177404
rect 220136 177364 262312 177392
rect 220136 177352 220142 177364
rect 262306 177352 262312 177364
rect 262364 177352 262370 177404
rect 289722 177352 289728 177404
rect 289780 177392 289786 177404
rect 310514 177392 310520 177404
rect 289780 177364 310520 177392
rect 289780 177352 289786 177364
rect 310514 177352 310520 177364
rect 310572 177352 310578 177404
rect 313918 177352 313924 177404
rect 313976 177392 313982 177404
rect 335538 177392 335544 177404
rect 313976 177364 335544 177392
rect 313976 177352 313982 177364
rect 335538 177352 335544 177364
rect 335596 177352 335602 177404
rect 166810 177284 166816 177336
rect 166868 177324 166874 177336
rect 197998 177324 198004 177336
rect 166868 177296 198004 177324
rect 166868 177284 166874 177296
rect 197998 177284 198004 177296
rect 198056 177284 198062 177336
rect 198182 177284 198188 177336
rect 198240 177324 198246 177336
rect 263594 177324 263600 177336
rect 198240 177296 263600 177324
rect 198240 177284 198246 177296
rect 263594 177284 263600 177296
rect 263652 177284 263658 177336
rect 287790 177284 287796 177336
rect 287848 177324 287854 177336
rect 334158 177324 334164 177336
rect 287848 177296 334164 177324
rect 287848 177284 287854 177296
rect 334158 177284 334164 177296
rect 334216 177284 334222 177336
rect 134426 177012 134432 177064
rect 134484 177052 134490 177064
rect 165246 177052 165252 177064
rect 134484 177024 165252 177052
rect 134484 177012 134490 177024
rect 165246 177012 165252 177024
rect 165304 177012 165310 177064
rect 127066 176944 127072 176996
rect 127124 176984 127130 176996
rect 173158 176984 173164 176996
rect 127124 176956 173164 176984
rect 127124 176944 127130 176956
rect 173158 176944 173164 176956
rect 173216 176944 173222 176996
rect 125778 176876 125784 176928
rect 125836 176916 125842 176928
rect 188338 176916 188344 176928
rect 125836 176888 188344 176916
rect 125836 176876 125842 176888
rect 188338 176876 188344 176888
rect 188396 176876 188402 176928
rect 108114 176808 108120 176860
rect 108172 176848 108178 176860
rect 170490 176848 170496 176860
rect 108172 176820 170496 176848
rect 108172 176808 108178 176820
rect 170490 176808 170496 176820
rect 170548 176808 170554 176860
rect 107010 176740 107016 176792
rect 107068 176780 107074 176792
rect 169294 176780 169300 176792
rect 107068 176752 169300 176780
rect 107068 176740 107074 176752
rect 169294 176740 169300 176752
rect 169352 176740 169358 176792
rect 135714 176672 135720 176724
rect 135772 176712 135778 176724
rect 135772 176684 212488 176712
rect 135772 176672 135778 176684
rect 212460 176644 212488 176684
rect 213914 176644 213920 176656
rect 212460 176616 213920 176644
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 235258 176604 235264 176656
rect 235316 176644 235322 176656
rect 248046 176644 248052 176656
rect 235316 176616 248052 176644
rect 235316 176604 235322 176616
rect 248046 176604 248052 176616
rect 248104 176604 248110 176656
rect 313826 176604 313832 176656
rect 313884 176644 313890 176656
rect 321462 176644 321468 176656
rect 313884 176616 321468 176644
rect 313884 176604 313890 176616
rect 321462 176604 321468 176616
rect 321520 176604 321526 176656
rect 319530 176536 319536 176588
rect 319588 176576 319594 176588
rect 321738 176576 321744 176588
rect 319588 176548 321744 176576
rect 319588 176536 319594 176548
rect 321738 176536 321744 176548
rect 321796 176536 321802 176588
rect 129458 176264 129464 176316
rect 129516 176304 129522 176316
rect 166166 176304 166172 176316
rect 129516 176276 166172 176304
rect 129516 176264 129522 176276
rect 166166 176264 166172 176276
rect 166224 176264 166230 176316
rect 119430 176196 119436 176248
rect 119488 176236 119494 176248
rect 166442 176236 166448 176248
rect 119488 176208 166448 176236
rect 119488 176196 119494 176208
rect 166442 176196 166448 176208
rect 166500 176196 166506 176248
rect 115750 176128 115756 176180
rect 115808 176168 115814 176180
rect 166258 176168 166264 176180
rect 115808 176140 166264 176168
rect 115808 176128 115814 176140
rect 166258 176128 166264 176140
rect 166316 176128 166322 176180
rect 98362 176060 98368 176112
rect 98420 176100 98426 176112
rect 169018 176100 169024 176112
rect 98420 176072 169024 176100
rect 98420 176060 98426 176072
rect 169018 176060 169024 176072
rect 169076 176060 169082 176112
rect 100754 175992 100760 176044
rect 100812 176032 100818 176044
rect 171870 176032 171876 176044
rect 100812 176004 171876 176032
rect 100812 175992 100818 176004
rect 171870 175992 171876 176004
rect 171928 175992 171934 176044
rect 13078 175924 13084 175976
rect 13136 175964 13142 175976
rect 111058 175964 111064 175976
rect 13136 175936 111064 175964
rect 13136 175924 13142 175936
rect 111058 175924 111064 175936
rect 111116 175924 111122 175976
rect 116946 175924 116952 175976
rect 117004 175964 117010 175976
rect 169110 175964 169116 175976
rect 117004 175936 169116 175964
rect 117004 175924 117010 175936
rect 169110 175924 169116 175936
rect 169168 175924 169174 175976
rect 246298 175924 246304 175976
rect 246356 175964 246362 175976
rect 252738 175964 252744 175976
rect 246356 175936 252744 175964
rect 246356 175924 246362 175936
rect 252738 175924 252744 175936
rect 252796 175924 252802 175976
rect 315390 175924 315396 175976
rect 315448 175964 315454 175976
rect 332870 175964 332876 175976
rect 315448 175936 332876 175964
rect 315448 175924 315454 175936
rect 332870 175924 332876 175936
rect 332928 175924 332934 175976
rect 166534 175244 166540 175296
rect 166592 175284 166598 175296
rect 343818 175284 343824 175296
rect 166592 175256 343824 175284
rect 166592 175244 166598 175256
rect 343818 175244 343824 175256
rect 343876 175244 343882 175296
rect 165246 175176 165252 175228
rect 165304 175216 165310 175228
rect 213914 175216 213920 175228
rect 165304 175188 213920 175216
rect 165304 175176 165310 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 164326 175108 164332 175160
rect 164384 175148 164390 175160
rect 214006 175148 214012 175160
rect 164384 175120 214012 175148
rect 164384 175108 164390 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 2774 164092 2780 164144
rect 2832 164132 2838 164144
rect 4798 164132 4804 164144
rect 2832 164104 4804 164132
rect 2832 164092 2838 164104
rect 4798 164092 4804 164104
rect 4856 164092 4862 164144
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 17218 150396 17224 150408
rect 3476 150368 17224 150396
rect 3476 150356 3482 150368
rect 17218 150356 17224 150368
rect 17276 150356 17282 150408
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 14458 137952 14464 137964
rect 3292 137924 14464 137952
rect 3292 137912 3298 137924
rect 14458 137912 14464 137924
rect 14516 137912 14522 137964
rect 63402 125604 63408 125656
rect 63460 125644 63466 125656
rect 66162 125644 66168 125656
rect 63460 125616 66168 125644
rect 63460 125604 63466 125616
rect 66162 125604 66168 125616
rect 66220 125604 66226 125656
rect 63310 121456 63316 121508
rect 63368 121496 63374 121508
rect 66070 121496 66076 121508
rect 63368 121468 66076 121496
rect 63368 121456 63374 121468
rect 66070 121456 66076 121468
rect 66128 121456 66134 121508
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 13078 111772 13084 111784
rect 3476 111744 13084 111772
rect 3476 111732 3482 111744
rect 13078 111732 13084 111744
rect 13136 111732 13142 111784
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 25498 97968 25504 97980
rect 3476 97940 25504 97968
rect 3476 97928 3482 97940
rect 25498 97928 25504 97940
rect 25556 97928 25562 97980
rect 262858 174496 262864 174548
rect 262916 174536 262922 174548
rect 274082 174536 274088 174548
rect 262916 174508 274088 174536
rect 262916 174496 262922 174508
rect 274082 174496 274088 174508
rect 274140 174496 274146 174548
rect 287974 174020 287980 174072
rect 288032 174060 288038 174072
rect 307570 174060 307576 174072
rect 288032 174032 307576 174060
rect 288032 174020 288038 174032
rect 307570 174020 307576 174032
rect 307628 174020 307634 174072
rect 271138 173952 271144 174004
rect 271196 173992 271202 174004
rect 307294 173992 307300 174004
rect 271196 173964 307300 173992
rect 271196 173952 271202 173964
rect 307294 173952 307300 173964
rect 307352 173952 307358 174004
rect 265894 173884 265900 173936
rect 265952 173924 265958 173936
rect 307662 173924 307668 173936
rect 265952 173896 307668 173924
rect 265952 173884 265958 173896
rect 307662 173884 307668 173896
rect 307720 173884 307726 173936
rect 165522 173816 165528 173868
rect 165580 173856 165586 173868
rect 214006 173856 214012 173868
rect 165580 173828 214012 173856
rect 165580 173816 165586 173828
rect 214006 173816 214012 173828
rect 214064 173816 214070 173868
rect 252462 173816 252468 173868
rect 252520 173856 252526 173868
rect 258074 173856 258080 173868
rect 252520 173828 258080 173856
rect 252520 173816 252526 173828
rect 258074 173816 258080 173828
rect 258132 173816 258138 173868
rect 167914 173748 167920 173800
rect 167972 173788 167978 173800
rect 213914 173788 213920 173800
rect 167972 173760 213920 173788
rect 167972 173748 167978 173760
rect 213914 173748 213920 173760
rect 213972 173748 213978 173800
rect 258074 173680 258080 173732
rect 258132 173720 258138 173732
rect 258350 173720 258356 173732
rect 258132 173692 258356 173720
rect 258132 173680 258138 173692
rect 258350 173680 258356 173692
rect 258408 173680 258414 173732
rect 251726 172796 251732 172848
rect 251784 172836 251790 172848
rect 255590 172836 255596 172848
rect 251784 172808 255596 172836
rect 251784 172796 251790 172808
rect 255590 172796 255596 172808
rect 255648 172796 255654 172848
rect 283650 172660 283656 172712
rect 283708 172700 283714 172712
rect 307570 172700 307576 172712
rect 283708 172672 307576 172700
rect 283708 172660 283714 172672
rect 307570 172660 307576 172672
rect 307628 172660 307634 172712
rect 269758 172592 269764 172644
rect 269816 172632 269822 172644
rect 307294 172632 307300 172644
rect 269816 172604 307300 172632
rect 269816 172592 269822 172604
rect 307294 172592 307300 172604
rect 307352 172592 307358 172644
rect 265710 172524 265716 172576
rect 265768 172564 265774 172576
rect 307662 172564 307668 172576
rect 265768 172536 307668 172564
rect 265768 172524 265774 172536
rect 307662 172524 307668 172536
rect 307720 172524 307726 172576
rect 166166 172456 166172 172508
rect 166224 172496 166230 172508
rect 213914 172496 213920 172508
rect 166224 172468 213920 172496
rect 166224 172456 166230 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 252462 172388 252468 172440
rect 252520 172428 252526 172440
rect 260834 172428 260840 172440
rect 252520 172400 260840 172428
rect 252520 172388 252526 172400
rect 260834 172388 260840 172400
rect 260892 172388 260898 172440
rect 252370 172320 252376 172372
rect 252428 172360 252434 172372
rect 262398 172360 262404 172372
rect 252428 172332 262404 172360
rect 252428 172320 252434 172332
rect 262398 172320 262404 172332
rect 262456 172320 262462 172372
rect 281074 171164 281080 171216
rect 281132 171204 281138 171216
rect 306926 171204 306932 171216
rect 281132 171176 306932 171204
rect 281132 171164 281138 171176
rect 306926 171164 306932 171176
rect 306984 171164 306990 171216
rect 262950 171096 262956 171148
rect 263008 171136 263014 171148
rect 307478 171136 307484 171148
rect 263008 171108 307484 171136
rect 263008 171096 263014 171108
rect 307478 171096 307484 171108
rect 307536 171096 307542 171148
rect 173158 171028 173164 171080
rect 173216 171068 173222 171080
rect 213914 171068 213920 171080
rect 173216 171040 213920 171068
rect 173216 171028 173222 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 188338 170960 188344 171012
rect 188396 171000 188402 171012
rect 214006 171000 214012 171012
rect 188396 170972 214012 171000
rect 188396 170960 188402 170972
rect 214006 170960 214012 170972
rect 214064 170960 214070 171012
rect 324314 170892 324320 170944
rect 324372 170932 324378 170944
rect 325970 170932 325976 170944
rect 324372 170904 325976 170932
rect 324372 170892 324378 170904
rect 325970 170892 325976 170904
rect 326028 170892 326034 170944
rect 251542 170756 251548 170808
rect 251600 170796 251606 170808
rect 254210 170796 254216 170808
rect 251600 170768 254216 170796
rect 251600 170756 251606 170768
rect 254210 170756 254216 170768
rect 254268 170756 254274 170808
rect 169294 170348 169300 170400
rect 169352 170388 169358 170400
rect 214834 170388 214840 170400
rect 169352 170360 214840 170388
rect 169352 170348 169358 170360
rect 214834 170348 214840 170360
rect 214892 170348 214898 170400
rect 252278 170280 252284 170332
rect 252336 170320 252342 170332
rect 256786 170320 256792 170332
rect 252336 170292 256792 170320
rect 252336 170280 252342 170292
rect 256786 170280 256792 170292
rect 256844 170280 256850 170332
rect 304258 169872 304264 169924
rect 304316 169912 304322 169924
rect 307478 169912 307484 169924
rect 304316 169884 307484 169912
rect 304316 169872 304322 169884
rect 307478 169872 307484 169884
rect 307536 169872 307542 169924
rect 273898 169804 273904 169856
rect 273956 169844 273962 169856
rect 307294 169844 307300 169856
rect 273956 169816 307300 169844
rect 273956 169804 273962 169816
rect 307294 169804 307300 169816
rect 307352 169804 307358 169856
rect 267182 169736 267188 169788
rect 267240 169776 267246 169788
rect 307662 169776 307668 169788
rect 267240 169748 307668 169776
rect 267240 169736 267246 169748
rect 307662 169736 307668 169748
rect 307720 169736 307726 169788
rect 166350 169668 166356 169720
rect 166408 169708 166414 169720
rect 213914 169708 213920 169720
rect 166408 169680 213920 169708
rect 166408 169668 166414 169680
rect 213914 169668 213920 169680
rect 213972 169668 213978 169720
rect 324314 169668 324320 169720
rect 324372 169708 324378 169720
rect 331214 169708 331220 169720
rect 324372 169680 331220 169708
rect 324372 169668 324378 169680
rect 331214 169668 331220 169680
rect 331272 169668 331278 169720
rect 252186 169600 252192 169652
rect 252244 169640 252250 169652
rect 258074 169640 258080 169652
rect 252244 169612 258080 169640
rect 252244 169600 252250 169612
rect 258074 169600 258080 169612
rect 258132 169600 258138 169652
rect 170490 168988 170496 169040
rect 170548 169028 170554 169040
rect 215018 169028 215024 169040
rect 170548 169000 215024 169028
rect 170548 168988 170554 169000
rect 215018 168988 215024 169000
rect 215076 168988 215082 169040
rect 287882 168512 287888 168564
rect 287940 168552 287946 168564
rect 307662 168552 307668 168564
rect 287940 168524 307668 168552
rect 287940 168512 287946 168524
rect 307662 168512 307668 168524
rect 307720 168512 307726 168564
rect 279418 168444 279424 168496
rect 279476 168484 279482 168496
rect 307570 168484 307576 168496
rect 279476 168456 307576 168484
rect 279476 168444 279482 168456
rect 307570 168444 307576 168456
rect 307628 168444 307634 168496
rect 264330 168376 264336 168428
rect 264388 168416 264394 168428
rect 307294 168416 307300 168428
rect 264388 168388 307300 168416
rect 264388 168376 264394 168388
rect 307294 168376 307300 168388
rect 307352 168376 307358 168428
rect 167730 168308 167736 168360
rect 167788 168348 167794 168360
rect 213914 168348 213920 168360
rect 167788 168320 213920 168348
rect 167788 168308 167794 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 252462 168308 252468 168360
rect 252520 168348 252526 168360
rect 263686 168348 263692 168360
rect 252520 168320 263692 168348
rect 252520 168308 252526 168320
rect 263686 168308 263692 168320
rect 263744 168308 263750 168360
rect 324314 168308 324320 168360
rect 324372 168348 324378 168360
rect 338390 168348 338396 168360
rect 324372 168320 338396 168348
rect 324372 168308 324378 168320
rect 338390 168308 338396 168320
rect 338448 168308 338454 168360
rect 211982 168240 211988 168292
rect 212040 168280 212046 168292
rect 214006 168280 214012 168292
rect 212040 168252 214012 168280
rect 212040 168240 212046 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 294598 167696 294604 167748
rect 294656 167736 294662 167748
rect 307018 167736 307024 167748
rect 294656 167708 307024 167736
rect 294656 167696 294662 167708
rect 307018 167696 307024 167708
rect 307076 167696 307082 167748
rect 258902 167628 258908 167680
rect 258960 167668 258966 167680
rect 307386 167668 307392 167680
rect 258960 167640 307392 167668
rect 258960 167628 258966 167640
rect 307386 167628 307392 167640
rect 307444 167628 307450 167680
rect 252278 167424 252284 167476
rect 252336 167464 252342 167476
rect 256694 167464 256700 167476
rect 252336 167436 256700 167464
rect 252336 167424 252342 167436
rect 256694 167424 256700 167436
rect 256752 167424 256758 167476
rect 267090 167016 267096 167068
rect 267148 167056 267154 167068
rect 306926 167056 306932 167068
rect 267148 167028 306932 167056
rect 267148 167016 267154 167028
rect 306926 167016 306932 167028
rect 306984 167016 306990 167068
rect 166442 166948 166448 167000
rect 166500 166988 166506 167000
rect 213914 166988 213920 167000
rect 166500 166960 213920 166988
rect 166500 166948 166506 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 167822 166880 167828 166932
rect 167880 166920 167886 166932
rect 214006 166920 214012 166932
rect 167880 166892 214012 166920
rect 167880 166880 167886 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 169110 166812 169116 166864
rect 169168 166852 169174 166864
rect 213914 166852 213920 166864
rect 169168 166824 213920 166852
rect 169168 166812 169174 166824
rect 213914 166812 213920 166824
rect 213972 166812 213978 166864
rect 252278 166812 252284 166864
rect 252336 166852 252342 166864
rect 258166 166852 258172 166864
rect 252336 166824 258172 166852
rect 252336 166812 252342 166824
rect 258166 166812 258172 166824
rect 258224 166812 258230 166864
rect 251910 166404 251916 166456
rect 251968 166444 251974 166456
rect 259546 166444 259552 166456
rect 251968 166416 259552 166444
rect 251968 166404 251974 166416
rect 259546 166404 259552 166416
rect 259604 166404 259610 166456
rect 249702 166268 249708 166320
rect 249760 166308 249766 166320
rect 305178 166308 305184 166320
rect 249760 166280 305184 166308
rect 249760 166268 249766 166280
rect 305178 166268 305184 166280
rect 305236 166268 305242 166320
rect 252278 166064 252284 166116
rect 252336 166104 252342 166116
rect 256878 166104 256884 166116
rect 252336 166076 256884 166104
rect 252336 166064 252342 166076
rect 256878 166064 256884 166076
rect 256936 166064 256942 166116
rect 282362 165724 282368 165776
rect 282420 165764 282426 165776
rect 306926 165764 306932 165776
rect 282420 165736 306932 165764
rect 282420 165724 282426 165736
rect 306926 165724 306932 165736
rect 306984 165724 306990 165776
rect 272518 165656 272524 165708
rect 272576 165696 272582 165708
rect 307478 165696 307484 165708
rect 272576 165668 307484 165696
rect 272576 165656 272582 165668
rect 307478 165656 307484 165668
rect 307536 165656 307542 165708
rect 257522 165588 257528 165640
rect 257580 165628 257586 165640
rect 307662 165628 307668 165640
rect 257580 165600 307668 165628
rect 257580 165588 257586 165600
rect 307662 165588 307668 165600
rect 307720 165588 307726 165640
rect 166258 165520 166264 165572
rect 166316 165560 166322 165572
rect 213914 165560 213920 165572
rect 166316 165532 213920 165560
rect 166316 165520 166322 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 252462 165520 252468 165572
rect 252520 165560 252526 165572
rect 270678 165560 270684 165572
rect 252520 165532 270684 165560
rect 252520 165520 252526 165532
rect 270678 165520 270684 165532
rect 270736 165520 270742 165572
rect 324406 165520 324412 165572
rect 324464 165560 324470 165572
rect 335354 165560 335360 165572
rect 324464 165532 335360 165560
rect 324464 165520 324470 165532
rect 335354 165520 335360 165532
rect 335412 165520 335418 165572
rect 209038 165452 209044 165504
rect 209096 165492 209102 165504
rect 214006 165492 214012 165504
rect 209096 165464 214012 165492
rect 209096 165452 209102 165464
rect 214006 165452 214012 165464
rect 214064 165452 214070 165504
rect 324314 165452 324320 165504
rect 324372 165492 324378 165504
rect 332870 165492 332876 165504
rect 324372 165464 332876 165492
rect 324372 165452 324378 165464
rect 332870 165452 332876 165464
rect 332928 165452 332934 165504
rect 251542 164432 251548 164484
rect 251600 164472 251606 164484
rect 252830 164472 252836 164484
rect 251600 164444 252836 164472
rect 251600 164432 251606 164444
rect 252830 164432 252836 164444
rect 252888 164432 252894 164484
rect 278130 164364 278136 164416
rect 278188 164404 278194 164416
rect 307662 164404 307668 164416
rect 278188 164376 307668 164404
rect 278188 164364 278194 164376
rect 307662 164364 307668 164376
rect 307720 164364 307726 164416
rect 271230 164296 271236 164348
rect 271288 164336 271294 164348
rect 307570 164336 307576 164348
rect 271288 164308 307576 164336
rect 271288 164296 271294 164308
rect 307570 164296 307576 164308
rect 307628 164296 307634 164348
rect 260190 164228 260196 164280
rect 260248 164268 260254 164280
rect 307294 164268 307300 164280
rect 260248 164240 307300 164268
rect 260248 164228 260254 164240
rect 307294 164228 307300 164240
rect 307352 164228 307358 164280
rect 211890 164160 211896 164212
rect 211948 164200 211954 164212
rect 213914 164200 213920 164212
rect 211948 164172 213920 164200
rect 211948 164160 211954 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 252462 164160 252468 164212
rect 252520 164200 252526 164212
rect 267826 164200 267832 164212
rect 252520 164172 267832 164200
rect 252520 164160 252526 164172
rect 267826 164160 267832 164172
rect 267884 164160 267890 164212
rect 324314 164160 324320 164212
rect 324372 164200 324378 164212
rect 339770 164200 339776 164212
rect 324372 164172 339776 164200
rect 324372 164160 324378 164172
rect 339770 164160 339776 164172
rect 339828 164160 339834 164212
rect 252094 164092 252100 164144
rect 252152 164132 252158 164144
rect 264974 164132 264980 164144
rect 252152 164104 264980 164132
rect 252152 164092 252158 164104
rect 264974 164092 264980 164104
rect 265032 164092 265038 164144
rect 324406 164092 324412 164144
rect 324464 164132 324470 164144
rect 334250 164132 334256 164144
rect 324464 164104 334256 164132
rect 324464 164092 324470 164104
rect 334250 164092 334256 164104
rect 334308 164092 334314 164144
rect 261110 163480 261116 163532
rect 261168 163520 261174 163532
rect 291838 163520 291844 163532
rect 261168 163492 291844 163520
rect 261168 163480 261174 163492
rect 291838 163480 291844 163492
rect 291896 163480 291902 163532
rect 290642 162936 290648 162988
rect 290700 162976 290706 162988
rect 307294 162976 307300 162988
rect 290700 162948 307300 162976
rect 290700 162936 290706 162948
rect 307294 162936 307300 162948
rect 307352 162936 307358 162988
rect 268470 162868 268476 162920
rect 268528 162908 268534 162920
rect 307662 162908 307668 162920
rect 268528 162880 307668 162908
rect 268528 162868 268534 162880
rect 307662 162868 307668 162880
rect 307720 162868 307726 162920
rect 252462 162800 252468 162852
rect 252520 162840 252526 162852
rect 270586 162840 270592 162852
rect 252520 162812 270592 162840
rect 252520 162800 252526 162812
rect 270586 162800 270592 162812
rect 270644 162800 270650 162852
rect 324314 162800 324320 162852
rect 324372 162840 324378 162852
rect 353294 162840 353300 162852
rect 324372 162812 353300 162840
rect 324372 162800 324378 162812
rect 353294 162800 353300 162812
rect 353352 162800 353358 162852
rect 263042 162120 263048 162172
rect 263100 162160 263106 162172
rect 307202 162160 307208 162172
rect 263100 162132 307208 162160
rect 263100 162120 263106 162132
rect 307202 162120 307208 162132
rect 307260 162120 307266 162172
rect 252462 161916 252468 161968
rect 252520 161956 252526 161968
rect 259638 161956 259644 161968
rect 252520 161928 259644 161956
rect 252520 161916 252526 161928
rect 259638 161916 259644 161928
rect 259696 161916 259702 161968
rect 298738 161508 298744 161560
rect 298796 161548 298802 161560
rect 307478 161548 307484 161560
rect 298796 161520 307484 161548
rect 298796 161508 298802 161520
rect 307478 161508 307484 161520
rect 307536 161508 307542 161560
rect 258810 161440 258816 161492
rect 258868 161480 258874 161492
rect 307662 161480 307668 161492
rect 258868 161452 307668 161480
rect 258868 161440 258874 161452
rect 307662 161440 307668 161452
rect 307720 161440 307726 161492
rect 324314 161372 324320 161424
rect 324372 161412 324378 161424
rect 341058 161412 341064 161424
rect 324372 161384 341064 161412
rect 324372 161372 324378 161384
rect 341058 161372 341064 161384
rect 341116 161372 341122 161424
rect 252462 161032 252468 161084
rect 252520 161072 252526 161084
rect 258258 161072 258264 161084
rect 252520 161044 258264 161072
rect 252520 161032 252526 161044
rect 258258 161032 258264 161044
rect 258316 161032 258322 161084
rect 252462 160896 252468 160948
rect 252520 160936 252526 160948
rect 259730 160936 259736 160948
rect 252520 160908 259736 160936
rect 252520 160896 252526 160908
rect 259730 160896 259736 160908
rect 259788 160896 259794 160948
rect 167914 160760 167920 160812
rect 167972 160800 167978 160812
rect 192662 160800 192668 160812
rect 167972 160772 192668 160800
rect 167972 160760 167978 160772
rect 192662 160760 192668 160772
rect 192720 160760 192726 160812
rect 177758 160692 177764 160744
rect 177816 160732 177822 160744
rect 215938 160732 215944 160744
rect 177816 160704 215944 160732
rect 177816 160692 177822 160704
rect 215938 160692 215944 160704
rect 215996 160692 216002 160744
rect 261478 160692 261484 160744
rect 261536 160732 261542 160744
rect 307110 160732 307116 160744
rect 261536 160704 307116 160732
rect 261536 160692 261542 160704
rect 307110 160692 307116 160704
rect 307168 160692 307174 160744
rect 302970 160216 302976 160268
rect 303028 160256 303034 160268
rect 307662 160256 307668 160268
rect 303028 160228 307668 160256
rect 303028 160216 303034 160228
rect 307662 160216 307668 160228
rect 307720 160216 307726 160268
rect 283742 160148 283748 160200
rect 283800 160188 283806 160200
rect 306742 160188 306748 160200
rect 283800 160160 306748 160188
rect 283800 160148 283806 160160
rect 306742 160148 306748 160160
rect 306800 160148 306806 160200
rect 253566 160080 253572 160132
rect 253624 160120 253630 160132
rect 255314 160120 255320 160132
rect 253624 160092 255320 160120
rect 253624 160080 253630 160092
rect 255314 160080 255320 160092
rect 255372 160080 255378 160132
rect 260098 160080 260104 160132
rect 260156 160120 260162 160132
rect 307478 160120 307484 160132
rect 260156 160092 307484 160120
rect 260156 160080 260162 160092
rect 307478 160080 307484 160092
rect 307536 160080 307542 160132
rect 169202 160012 169208 160064
rect 169260 160052 169266 160064
rect 213914 160052 213920 160064
rect 169260 160024 213920 160052
rect 169260 160012 169266 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 252462 160012 252468 160064
rect 252520 160052 252526 160064
rect 269206 160052 269212 160064
rect 252520 160024 269212 160052
rect 252520 160012 252526 160024
rect 269206 160012 269212 160024
rect 269264 160012 269270 160064
rect 324314 160012 324320 160064
rect 324372 160052 324378 160064
rect 331398 160052 331404 160064
rect 324372 160024 331404 160052
rect 324372 160012 324378 160024
rect 331398 160012 331404 160024
rect 331456 160012 331462 160064
rect 173250 159944 173256 159996
rect 173308 159984 173314 159996
rect 214006 159984 214012 159996
rect 173308 159956 214012 159984
rect 173308 159944 173314 159956
rect 214006 159944 214012 159956
rect 214064 159944 214070 159996
rect 251910 159944 251916 159996
rect 251968 159984 251974 159996
rect 266446 159984 266452 159996
rect 251968 159956 266452 159984
rect 251968 159944 251974 159956
rect 266446 159944 266452 159956
rect 266504 159944 266510 159996
rect 258994 159332 259000 159384
rect 259052 159372 259058 159384
rect 307386 159372 307392 159384
rect 259052 159344 307392 159372
rect 259052 159332 259058 159344
rect 307386 159332 307392 159344
rect 307444 159332 307450 159384
rect 301498 158788 301504 158840
rect 301556 158828 301562 158840
rect 307662 158828 307668 158840
rect 301556 158800 307668 158828
rect 301556 158788 301562 158800
rect 307662 158788 307668 158800
rect 307720 158788 307726 158840
rect 265802 158720 265808 158772
rect 265860 158760 265866 158772
rect 307570 158760 307576 158772
rect 265860 158732 307576 158760
rect 265860 158720 265866 158732
rect 307570 158720 307576 158732
rect 307628 158720 307634 158772
rect 184198 158652 184204 158704
rect 184256 158692 184262 158704
rect 213914 158692 213920 158704
rect 184256 158664 213920 158692
rect 184256 158652 184262 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 324406 158652 324412 158704
rect 324464 158692 324470 158704
rect 343910 158692 343916 158704
rect 324464 158664 343916 158692
rect 324464 158652 324470 158664
rect 343910 158652 343916 158664
rect 343968 158652 343974 158704
rect 324314 158584 324320 158636
rect 324372 158624 324378 158636
rect 332778 158624 332784 158636
rect 324372 158596 332784 158624
rect 324372 158584 324378 158596
rect 332778 158584 332784 158596
rect 332836 158584 332842 158636
rect 252554 157972 252560 158024
rect 252612 158012 252618 158024
rect 260926 158012 260932 158024
rect 252612 157984 260932 158012
rect 252612 157972 252618 157984
rect 260926 157972 260932 157984
rect 260984 157972 260990 158024
rect 296070 157496 296076 157548
rect 296128 157536 296134 157548
rect 307662 157536 307668 157548
rect 296128 157508 307668 157536
rect 296128 157496 296134 157508
rect 307662 157496 307668 157508
rect 307720 157496 307726 157548
rect 264422 157428 264428 157480
rect 264480 157468 264486 157480
rect 306926 157468 306932 157480
rect 264480 157440 306932 157468
rect 264480 157428 264486 157440
rect 306926 157428 306932 157440
rect 306984 157428 306990 157480
rect 257430 157360 257436 157412
rect 257488 157400 257494 157412
rect 307294 157400 307300 157412
rect 257488 157372 307300 157400
rect 257488 157360 257494 157372
rect 307294 157360 307300 157372
rect 307352 157360 307358 157412
rect 170398 157292 170404 157344
rect 170456 157332 170462 157344
rect 214006 157332 214012 157344
rect 170456 157304 214012 157332
rect 170456 157292 170462 157304
rect 214006 157292 214012 157304
rect 214064 157292 214070 157344
rect 251542 157292 251548 157344
rect 251600 157332 251606 157344
rect 274818 157332 274824 157344
rect 251600 157304 274824 157332
rect 251600 157292 251606 157304
rect 274818 157292 274824 157304
rect 274876 157292 274882 157344
rect 324314 157292 324320 157344
rect 324372 157332 324378 157344
rect 336918 157332 336924 157344
rect 324372 157304 336924 157332
rect 324372 157292 324378 157304
rect 336918 157292 336924 157304
rect 336976 157292 336982 157344
rect 171870 157224 171876 157276
rect 171928 157264 171934 157276
rect 213914 157264 213920 157276
rect 171928 157236 213920 157264
rect 171928 157224 171934 157236
rect 213914 157224 213920 157236
rect 213972 157224 213978 157276
rect 252462 157224 252468 157276
rect 252520 157264 252526 157276
rect 269298 157264 269304 157276
rect 252520 157236 269304 157264
rect 252520 157224 252526 157236
rect 269298 157224 269304 157236
rect 269356 157224 269362 157276
rect 324406 157156 324412 157208
rect 324464 157196 324470 157208
rect 327350 157196 327356 157208
rect 324464 157168 327356 157196
rect 324464 157156 324470 157168
rect 327350 157156 327356 157168
rect 327408 157156 327414 157208
rect 278406 156612 278412 156664
rect 278464 156652 278470 156664
rect 307662 156652 307668 156664
rect 278464 156624 307668 156652
rect 278464 156612 278470 156624
rect 307662 156612 307668 156624
rect 307720 156612 307726 156664
rect 269850 156000 269856 156052
rect 269908 156040 269914 156052
rect 307478 156040 307484 156052
rect 269908 156012 307484 156040
rect 269908 156000 269914 156012
rect 307478 156000 307484 156012
rect 307536 156000 307542 156052
rect 261570 155932 261576 155984
rect 261628 155972 261634 155984
rect 306742 155972 306748 155984
rect 261628 155944 306748 155972
rect 261628 155932 261634 155944
rect 306742 155932 306748 155944
rect 306800 155932 306806 155984
rect 169018 155864 169024 155916
rect 169076 155904 169082 155916
rect 213914 155904 213920 155916
rect 169076 155876 213920 155904
rect 169076 155864 169082 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 252370 155864 252376 155916
rect 252428 155904 252434 155916
rect 276106 155904 276112 155916
rect 252428 155876 276112 155904
rect 252428 155864 252434 155876
rect 276106 155864 276112 155876
rect 276164 155864 276170 155916
rect 324314 155864 324320 155916
rect 324372 155904 324378 155916
rect 356054 155904 356060 155916
rect 324372 155876 356060 155904
rect 324372 155864 324378 155876
rect 356054 155864 356060 155876
rect 356112 155864 356118 155916
rect 252462 155796 252468 155848
rect 252520 155836 252526 155848
rect 263594 155836 263600 155848
rect 252520 155808 263600 155836
rect 252520 155796 252526 155808
rect 263594 155796 263600 155808
rect 263652 155796 263658 155848
rect 204898 155184 204904 155236
rect 204956 155224 204962 155236
rect 216122 155224 216128 155236
rect 204956 155196 216128 155224
rect 204956 155184 204962 155196
rect 216122 155184 216128 155196
rect 216180 155184 216186 155236
rect 251726 155184 251732 155236
rect 251784 155224 251790 155236
rect 269114 155224 269120 155236
rect 251784 155196 269120 155224
rect 251784 155184 251790 155196
rect 269114 155184 269120 155196
rect 269172 155184 269178 155236
rect 285214 154708 285220 154760
rect 285272 154748 285278 154760
rect 307570 154748 307576 154760
rect 285272 154720 307576 154748
rect 285272 154708 285278 154720
rect 307570 154708 307576 154720
rect 307628 154708 307634 154760
rect 276750 154640 276756 154692
rect 276808 154680 276814 154692
rect 307662 154680 307668 154692
rect 276808 154652 307668 154680
rect 276808 154640 276814 154652
rect 307662 154640 307668 154652
rect 307720 154640 307726 154692
rect 253474 154572 253480 154624
rect 253532 154612 253538 154624
rect 307478 154612 307484 154624
rect 253532 154584 307484 154612
rect 253532 154572 253538 154584
rect 307478 154572 307484 154584
rect 307536 154572 307542 154624
rect 252002 154504 252008 154556
rect 252060 154544 252066 154556
rect 277394 154544 277400 154556
rect 252060 154516 277400 154544
rect 252060 154504 252066 154516
rect 277394 154504 277400 154516
rect 277452 154504 277458 154556
rect 324314 154504 324320 154556
rect 324372 154544 324378 154556
rect 346578 154544 346584 154556
rect 324372 154516 346584 154544
rect 324372 154504 324378 154516
rect 346578 154504 346584 154516
rect 346636 154504 346642 154556
rect 251542 154436 251548 154488
rect 251600 154476 251606 154488
rect 272058 154476 272064 154488
rect 251600 154448 272064 154476
rect 251600 154436 251606 154448
rect 272058 154436 272064 154448
rect 272116 154436 272122 154488
rect 324406 154436 324412 154488
rect 324464 154476 324470 154488
rect 330110 154476 330116 154488
rect 324464 154448 330116 154476
rect 324464 154436 324470 154448
rect 330110 154436 330116 154448
rect 330168 154436 330174 154488
rect 252462 154368 252468 154420
rect 252520 154408 252526 154420
rect 267918 154408 267924 154420
rect 252520 154380 267924 154408
rect 252520 154368 252526 154380
rect 267918 154368 267924 154380
rect 267976 154368 267982 154420
rect 282454 153824 282460 153876
rect 282512 153864 282518 153876
rect 307386 153864 307392 153876
rect 282512 153836 307392 153864
rect 282512 153824 282518 153836
rect 307386 153824 307392 153836
rect 307444 153824 307450 153876
rect 204990 153280 204996 153332
rect 205048 153320 205054 153332
rect 214006 153320 214012 153332
rect 205048 153292 214012 153320
rect 205048 153280 205054 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 269942 153280 269948 153332
rect 270000 153320 270006 153332
rect 307662 153320 307668 153332
rect 270000 153292 307668 153320
rect 270000 153280 270006 153292
rect 307662 153280 307668 153292
rect 307720 153280 307726 153332
rect 202138 153212 202144 153264
rect 202196 153252 202202 153264
rect 213914 153252 213920 153264
rect 202196 153224 213920 153252
rect 202196 153212 202202 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 261662 153212 261668 153264
rect 261720 153252 261726 153264
rect 307478 153252 307484 153264
rect 261720 153224 307484 153252
rect 261720 153212 261726 153224
rect 307478 153212 307484 153224
rect 307536 153212 307542 153264
rect 252278 153144 252284 153196
rect 252336 153184 252342 153196
rect 278958 153184 278964 153196
rect 252336 153156 278964 153184
rect 252336 153144 252342 153156
rect 278958 153144 278964 153156
rect 279016 153144 279022 153196
rect 324314 153144 324320 153196
rect 324372 153184 324378 153196
rect 341150 153184 341156 153196
rect 324372 153156 341156 153184
rect 324372 153144 324378 153156
rect 341150 153144 341156 153156
rect 341208 153144 341214 153196
rect 250806 152668 250812 152720
rect 250864 152708 250870 152720
rect 258350 152708 258356 152720
rect 250864 152680 258356 152708
rect 250864 152668 250870 152680
rect 258350 152668 258356 152680
rect 258408 152668 258414 152720
rect 250530 152600 250536 152652
rect 250588 152640 250594 152652
rect 261018 152640 261024 152652
rect 250588 152612 261024 152640
rect 250588 152600 250594 152612
rect 261018 152600 261024 152612
rect 261076 152600 261082 152652
rect 251818 152532 251824 152584
rect 251876 152572 251882 152584
rect 272518 152572 272524 152584
rect 251876 152544 272524 152572
rect 251876 152532 251882 152544
rect 272518 152532 272524 152544
rect 272576 152532 272582 152584
rect 255958 152464 255964 152516
rect 256016 152504 256022 152516
rect 307570 152504 307576 152516
rect 256016 152476 307576 152504
rect 256016 152464 256022 152476
rect 307570 152464 307576 152476
rect 307628 152464 307634 152516
rect 195238 151852 195244 151904
rect 195296 151892 195302 151904
rect 213914 151892 213920 151904
rect 195296 151864 213920 151892
rect 195296 151852 195302 151864
rect 213914 151852 213920 151864
rect 213972 151852 213978 151904
rect 285122 151852 285128 151904
rect 285180 151892 285186 151904
rect 307478 151892 307484 151904
rect 285180 151864 307484 151892
rect 285180 151852 285186 151864
rect 307478 151852 307484 151864
rect 307536 151852 307542 151904
rect 184198 151784 184204 151836
rect 184256 151824 184262 151836
rect 214006 151824 214012 151836
rect 184256 151796 214012 151824
rect 184256 151784 184262 151796
rect 214006 151784 214012 151796
rect 214064 151784 214070 151836
rect 275554 151784 275560 151836
rect 275612 151824 275618 151836
rect 307662 151824 307668 151836
rect 275612 151796 307668 151824
rect 275612 151784 275618 151796
rect 307662 151784 307668 151796
rect 307720 151784 307726 151836
rect 324406 151716 324412 151768
rect 324464 151756 324470 151768
rect 336826 151756 336832 151768
rect 324464 151728 336832 151756
rect 324464 151716 324470 151728
rect 336826 151716 336832 151728
rect 336884 151716 336890 151768
rect 252370 151648 252376 151700
rect 252428 151688 252434 151700
rect 262306 151688 262312 151700
rect 252428 151660 262312 151688
rect 252428 151648 252434 151660
rect 262306 151648 262312 151660
rect 262364 151648 262370 151700
rect 324314 151648 324320 151700
rect 324372 151688 324378 151700
rect 328638 151688 328644 151700
rect 324372 151660 328644 151688
rect 324372 151648 324378 151660
rect 328638 151648 328644 151660
rect 328696 151648 328702 151700
rect 252462 151580 252468 151632
rect 252520 151620 252526 151632
rect 273346 151620 273352 151632
rect 252520 151592 273352 151620
rect 252520 151580 252526 151592
rect 273346 151580 273352 151592
rect 273404 151580 273410 151632
rect 251266 151240 251272 151292
rect 251324 151280 251330 151292
rect 253934 151280 253940 151292
rect 251324 151252 253940 151280
rect 251324 151240 251330 151252
rect 253934 151240 253940 151252
rect 253992 151240 253998 151292
rect 177850 151036 177856 151088
rect 177908 151076 177914 151088
rect 211798 151076 211804 151088
rect 177908 151048 211804 151076
rect 177908 151036 177914 151048
rect 211798 151036 211804 151048
rect 211856 151036 211862 151088
rect 256326 151036 256332 151088
rect 256384 151076 256390 151088
rect 306650 151076 306656 151088
rect 256384 151048 306656 151076
rect 256384 151036 256390 151048
rect 306650 151036 306656 151048
rect 306708 151036 306714 151088
rect 274174 150492 274180 150544
rect 274232 150532 274238 150544
rect 307478 150532 307484 150544
rect 274232 150504 307484 150532
rect 274232 150492 274238 150504
rect 307478 150492 307484 150504
rect 307536 150492 307542 150544
rect 206370 150424 206376 150476
rect 206428 150464 206434 150476
rect 213914 150464 213920 150476
rect 206428 150436 213920 150464
rect 206428 150424 206434 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 258718 150424 258724 150476
rect 258776 150464 258782 150476
rect 307662 150464 307668 150476
rect 258776 150436 307668 150464
rect 258776 150424 258782 150436
rect 307662 150424 307668 150436
rect 307720 150424 307726 150476
rect 192662 150356 192668 150408
rect 192720 150396 192726 150408
rect 214006 150396 214012 150408
rect 192720 150368 214012 150396
rect 192720 150356 192726 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 252462 150356 252468 150408
rect 252520 150396 252526 150408
rect 274726 150396 274732 150408
rect 252520 150368 274732 150396
rect 252520 150356 252526 150368
rect 274726 150356 274732 150368
rect 274784 150356 274790 150408
rect 324314 150356 324320 150408
rect 324372 150396 324378 150408
rect 346670 150396 346676 150408
rect 324372 150368 346676 150396
rect 324372 150356 324378 150368
rect 346670 150356 346676 150368
rect 346728 150356 346734 150408
rect 254670 149676 254676 149728
rect 254728 149716 254734 149728
rect 306558 149716 306564 149728
rect 254728 149688 306564 149716
rect 254728 149676 254734 149688
rect 306558 149676 306564 149688
rect 306616 149676 306622 149728
rect 251726 149608 251732 149660
rect 251784 149648 251790 149660
rect 255498 149648 255504 149660
rect 251784 149620 255504 149648
rect 251784 149608 251790 149620
rect 255498 149608 255504 149620
rect 255556 149608 255562 149660
rect 303154 149200 303160 149252
rect 303212 149240 303218 149252
rect 307294 149240 307300 149252
rect 303212 149212 307300 149240
rect 303212 149200 303218 149212
rect 307294 149200 307300 149212
rect 307352 149200 307358 149252
rect 276658 149132 276664 149184
rect 276716 149172 276722 149184
rect 306926 149172 306932 149184
rect 276716 149144 306932 149172
rect 276716 149132 276722 149144
rect 306926 149132 306932 149144
rect 306984 149132 306990 149184
rect 260374 149064 260380 149116
rect 260432 149104 260438 149116
rect 307478 149104 307484 149116
rect 260432 149076 307484 149104
rect 260432 149064 260438 149076
rect 307478 149064 307484 149076
rect 307536 149064 307542 149116
rect 167638 148996 167644 149048
rect 167696 149036 167702 149048
rect 213914 149036 213920 149048
rect 167696 149008 213920 149036
rect 167696 148996 167702 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 252462 148996 252468 149048
rect 252520 149036 252526 149048
rect 280154 149036 280160 149048
rect 252520 149008 280160 149036
rect 252520 148996 252526 149008
rect 280154 148996 280160 149008
rect 280212 148996 280218 149048
rect 324314 148996 324320 149048
rect 324372 149036 324378 149048
rect 338298 149036 338304 149048
rect 324372 149008 338304 149036
rect 324372 148996 324378 149008
rect 338298 148996 338304 149008
rect 338356 148996 338362 149048
rect 251542 148384 251548 148436
rect 251600 148424 251606 148436
rect 255406 148424 255412 148436
rect 251600 148396 255412 148424
rect 251600 148384 251606 148396
rect 255406 148384 255412 148396
rect 255464 148384 255470 148436
rect 254762 148316 254768 148368
rect 254820 148356 254826 148368
rect 307202 148356 307208 148368
rect 254820 148328 307208 148356
rect 254820 148316 254826 148328
rect 307202 148316 307208 148328
rect 307260 148316 307266 148368
rect 252370 147704 252376 147756
rect 252428 147744 252434 147756
rect 256970 147744 256976 147756
rect 252428 147716 256976 147744
rect 252428 147704 252434 147716
rect 256970 147704 256976 147716
rect 257028 147704 257034 147756
rect 272610 147704 272616 147756
rect 272668 147744 272674 147756
rect 307478 147744 307484 147756
rect 272668 147716 307484 147744
rect 272668 147704 272674 147716
rect 307478 147704 307484 147716
rect 307536 147704 307542 147756
rect 185670 147636 185676 147688
rect 185728 147676 185734 147688
rect 213914 147676 213920 147688
rect 185728 147648 213920 147676
rect 185728 147636 185734 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 257338 147636 257344 147688
rect 257396 147676 257402 147688
rect 307662 147676 307668 147688
rect 257396 147648 307668 147676
rect 257396 147636 257402 147648
rect 307662 147636 307668 147648
rect 307720 147636 307726 147688
rect 252462 147568 252468 147620
rect 252520 147608 252526 147620
rect 267734 147608 267740 147620
rect 252520 147580 267740 147608
rect 252520 147568 252526 147580
rect 267734 147568 267740 147580
rect 267792 147568 267798 147620
rect 324314 147568 324320 147620
rect 324372 147608 324378 147620
rect 347774 147608 347780 147620
rect 324372 147580 347780 147608
rect 324372 147568 324378 147580
rect 347774 147568 347780 147580
rect 347832 147568 347838 147620
rect 251266 147228 251272 147280
rect 251324 147268 251330 147280
rect 254026 147268 254032 147280
rect 251324 147240 254032 147268
rect 251324 147228 251330 147240
rect 254026 147228 254032 147240
rect 254084 147228 254090 147280
rect 177298 146888 177304 146940
rect 177356 146928 177362 146940
rect 214098 146928 214104 146940
rect 177356 146900 214104 146928
rect 177356 146888 177362 146900
rect 214098 146888 214104 146900
rect 214156 146888 214162 146940
rect 284938 146412 284944 146464
rect 284996 146452 285002 146464
rect 307662 146452 307668 146464
rect 284996 146424 307668 146452
rect 284996 146412 285002 146424
rect 307662 146412 307668 146424
rect 307720 146412 307726 146464
rect 256234 146344 256240 146396
rect 256292 146384 256298 146396
rect 306742 146384 306748 146396
rect 256292 146356 306748 146384
rect 256292 146344 256298 146356
rect 306742 146344 306748 146356
rect 306800 146344 306806 146396
rect 203518 146276 203524 146328
rect 203576 146316 203582 146328
rect 213914 146316 213920 146328
rect 203576 146288 213920 146316
rect 203576 146276 203582 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 256142 146276 256148 146328
rect 256200 146316 256206 146328
rect 307570 146316 307576 146328
rect 256200 146288 307576 146316
rect 256200 146276 256206 146288
rect 307570 146276 307576 146288
rect 307628 146276 307634 146328
rect 252462 146208 252468 146260
rect 252520 146248 252526 146260
rect 276014 146248 276020 146260
rect 252520 146220 276020 146248
rect 252520 146208 252526 146220
rect 276014 146208 276020 146220
rect 276072 146208 276078 146260
rect 252094 146140 252100 146192
rect 252152 146180 252158 146192
rect 273254 146180 273260 146192
rect 252152 146152 273260 146180
rect 252152 146140 252158 146152
rect 273254 146140 273260 146152
rect 273312 146140 273318 146192
rect 261754 145528 261760 145580
rect 261812 145568 261818 145580
rect 307018 145568 307024 145580
rect 261812 145540 307024 145568
rect 261812 145528 261818 145540
rect 307018 145528 307024 145540
rect 307076 145528 307082 145580
rect 211890 144984 211896 145036
rect 211948 145024 211954 145036
rect 214466 145024 214472 145036
rect 211948 144996 214472 145024
rect 211948 144984 211954 144996
rect 214466 144984 214472 144996
rect 214524 144984 214530 145036
rect 299014 144984 299020 145036
rect 299072 145024 299078 145036
rect 307478 145024 307484 145036
rect 299072 144996 307484 145024
rect 299072 144984 299078 144996
rect 307478 144984 307484 144996
rect 307536 144984 307542 145036
rect 170398 144916 170404 144968
rect 170456 144956 170462 144968
rect 213914 144956 213920 144968
rect 170456 144928 213920 144956
rect 170456 144916 170462 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 254578 144916 254584 144968
rect 254636 144956 254642 144968
rect 307662 144956 307668 144968
rect 254636 144928 307668 144956
rect 254636 144916 254642 144928
rect 307662 144916 307668 144928
rect 307720 144916 307726 144968
rect 252462 144848 252468 144900
rect 252520 144888 252526 144900
rect 266354 144888 266360 144900
rect 252520 144860 266360 144888
rect 252520 144848 252526 144860
rect 266354 144848 266360 144860
rect 266412 144848 266418 144900
rect 324314 144848 324320 144900
rect 324372 144888 324378 144900
rect 345198 144888 345204 144900
rect 324372 144860 345204 144888
rect 324372 144848 324378 144860
rect 345198 144848 345204 144860
rect 345256 144848 345262 144900
rect 252094 144780 252100 144832
rect 252152 144820 252158 144832
rect 262214 144820 262220 144832
rect 252152 144792 262220 144820
rect 252152 144780 252158 144792
rect 262214 144780 262220 144792
rect 262272 144780 262278 144832
rect 299106 144168 299112 144220
rect 299164 144208 299170 144220
rect 307294 144208 307300 144220
rect 299164 144180 307300 144208
rect 299164 144168 299170 144180
rect 307294 144168 307300 144180
rect 307352 144168 307358 144220
rect 251542 143624 251548 143676
rect 251600 143664 251606 143676
rect 259454 143664 259460 143676
rect 251600 143636 259460 143664
rect 251600 143624 251606 143636
rect 259454 143624 259460 143636
rect 259512 143624 259518 143676
rect 279602 143624 279608 143676
rect 279660 143664 279666 143676
rect 307478 143664 307484 143676
rect 279660 143636 307484 143664
rect 279660 143624 279666 143636
rect 307478 143624 307484 143636
rect 307536 143624 307542 143676
rect 167638 143556 167644 143608
rect 167696 143596 167702 143608
rect 213914 143596 213920 143608
rect 167696 143568 213920 143596
rect 167696 143556 167702 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 253382 143556 253388 143608
rect 253440 143596 253446 143608
rect 306926 143596 306932 143608
rect 253440 143568 306932 143596
rect 253440 143556 253446 143568
rect 306926 143556 306932 143568
rect 306984 143556 306990 143608
rect 324314 143488 324320 143540
rect 324372 143528 324378 143540
rect 335538 143528 335544 143540
rect 324372 143500 335544 143528
rect 324372 143488 324378 143500
rect 335538 143488 335544 143500
rect 335596 143488 335602 143540
rect 251910 142808 251916 142860
rect 251968 142848 251974 142860
rect 269850 142848 269856 142860
rect 251968 142820 269856 142848
rect 251968 142808 251974 142820
rect 269850 142808 269856 142820
rect 269908 142808 269914 142860
rect 301682 142264 301688 142316
rect 301740 142304 301746 142316
rect 307386 142304 307392 142316
rect 301740 142276 307392 142304
rect 301740 142264 301746 142276
rect 307386 142264 307392 142276
rect 307444 142264 307450 142316
rect 271322 142196 271328 142248
rect 271380 142236 271386 142248
rect 306742 142236 306748 142248
rect 271380 142208 306748 142236
rect 271380 142196 271386 142208
rect 306742 142196 306748 142208
rect 306800 142196 306806 142248
rect 209038 142128 209044 142180
rect 209096 142168 209102 142180
rect 213914 142168 213920 142180
rect 209096 142140 213920 142168
rect 209096 142128 209102 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 253290 142128 253296 142180
rect 253348 142168 253354 142180
rect 307662 142168 307668 142180
rect 253348 142140 307668 142168
rect 253348 142128 253354 142140
rect 307662 142128 307668 142140
rect 307720 142128 307726 142180
rect 252462 141924 252468 141976
rect 252520 141964 252526 141976
rect 256786 141964 256792 141976
rect 252520 141936 256792 141964
rect 252520 141924 252526 141936
rect 256786 141924 256792 141936
rect 256844 141924 256850 141976
rect 262858 141380 262864 141432
rect 262916 141420 262922 141432
rect 306558 141420 306564 141432
rect 262916 141392 306564 141420
rect 262916 141380 262922 141392
rect 306558 141380 306564 141392
rect 306616 141380 306622 141432
rect 304350 140904 304356 140956
rect 304408 140944 304414 140956
rect 307662 140944 307668 140956
rect 304408 140916 307668 140944
rect 304408 140904 304414 140916
rect 307662 140904 307668 140916
rect 307720 140904 307726 140956
rect 289354 140836 289360 140888
rect 289412 140876 289418 140888
rect 307570 140876 307576 140888
rect 289412 140848 307576 140876
rect 289412 140836 289418 140848
rect 307570 140836 307576 140848
rect 307628 140836 307634 140888
rect 182818 140768 182824 140820
rect 182876 140808 182882 140820
rect 213914 140808 213920 140820
rect 182876 140780 213920 140808
rect 182876 140768 182882 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 275462 140768 275468 140820
rect 275520 140808 275526 140820
rect 307478 140808 307484 140820
rect 275520 140780 307484 140808
rect 275520 140768 275526 140780
rect 307478 140768 307484 140780
rect 307536 140768 307542 140820
rect 251174 140428 251180 140480
rect 251232 140468 251238 140480
rect 253566 140468 253572 140480
rect 251232 140440 253572 140468
rect 251232 140428 251238 140440
rect 253566 140428 253572 140440
rect 253624 140428 253630 140480
rect 184474 140020 184480 140072
rect 184532 140060 184538 140072
rect 214650 140060 214656 140072
rect 184532 140032 214656 140060
rect 184532 140020 184538 140032
rect 214650 140020 214656 140032
rect 214708 140020 214714 140072
rect 193858 139476 193864 139528
rect 193916 139516 193922 139528
rect 214006 139516 214012 139528
rect 193916 139488 214012 139516
rect 193916 139476 193922 139488
rect 214006 139476 214012 139488
rect 214064 139476 214070 139528
rect 181438 139408 181444 139460
rect 181496 139448 181502 139460
rect 213914 139448 213920 139460
rect 181496 139420 213920 139448
rect 181496 139408 181502 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 280890 139408 280896 139460
rect 280948 139448 280954 139460
rect 307662 139448 307668 139460
rect 280948 139420 307668 139448
rect 280948 139408 280954 139420
rect 307662 139408 307668 139420
rect 307720 139408 307726 139460
rect 252462 139340 252468 139392
rect 252520 139380 252526 139392
rect 278866 139380 278872 139392
rect 252520 139352 278872 139380
rect 252520 139340 252526 139352
rect 278866 139340 278872 139352
rect 278924 139340 278930 139392
rect 324314 139340 324320 139392
rect 324372 139380 324378 139392
rect 338206 139380 338212 139392
rect 324372 139352 338212 139380
rect 324372 139340 324378 139352
rect 338206 139340 338212 139352
rect 338264 139340 338270 139392
rect 468478 139340 468484 139392
rect 468536 139380 468542 139392
rect 580166 139380 580172 139392
rect 468536 139352 580172 139380
rect 468536 139340 468542 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 251726 138728 251732 138780
rect 251784 138768 251790 138780
rect 271138 138768 271144 138780
rect 251784 138740 271144 138768
rect 251784 138728 251790 138740
rect 271138 138728 271144 138740
rect 271196 138728 271202 138780
rect 250714 138660 250720 138712
rect 250772 138700 250778 138712
rect 300946 138700 300952 138712
rect 250772 138672 300952 138700
rect 250772 138660 250778 138672
rect 300946 138660 300952 138672
rect 301004 138660 301010 138712
rect 297542 138116 297548 138168
rect 297600 138156 297606 138168
rect 307662 138156 307668 138168
rect 297600 138128 307668 138156
rect 297600 138116 297606 138128
rect 307662 138116 307668 138128
rect 307720 138116 307726 138168
rect 207658 138048 207664 138100
rect 207716 138088 207722 138100
rect 214006 138088 214012 138100
rect 207716 138060 214012 138088
rect 207716 138048 207722 138060
rect 214006 138048 214012 138060
rect 214064 138048 214070 138100
rect 290550 138048 290556 138100
rect 290608 138088 290614 138100
rect 307570 138088 307576 138100
rect 290608 138060 307576 138088
rect 290608 138048 290614 138060
rect 307570 138048 307576 138060
rect 307628 138048 307634 138100
rect 192662 137980 192668 138032
rect 192720 138020 192726 138032
rect 213914 138020 213920 138032
rect 192720 137992 213920 138020
rect 192720 137980 192726 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 272518 137980 272524 138032
rect 272576 138020 272582 138032
rect 307478 138020 307484 138032
rect 272576 137992 307484 138020
rect 272576 137980 272582 137992
rect 307478 137980 307484 137992
rect 307536 137980 307542 138032
rect 252462 137912 252468 137964
rect 252520 137952 252526 137964
rect 271966 137952 271972 137964
rect 252520 137924 271972 137952
rect 252520 137912 252526 137924
rect 271966 137912 271972 137924
rect 272024 137912 272030 137964
rect 324314 137912 324320 137964
rect 324372 137952 324378 137964
rect 345106 137952 345112 137964
rect 324372 137924 345112 137952
rect 324372 137912 324378 137924
rect 345106 137912 345112 137924
rect 345164 137912 345170 137964
rect 324498 137844 324504 137896
rect 324556 137884 324562 137896
rect 328546 137884 328552 137896
rect 324556 137856 328552 137884
rect 324556 137844 324562 137856
rect 328546 137844 328552 137856
rect 328604 137844 328610 137896
rect 251266 137708 251272 137760
rect 251324 137748 251330 137760
rect 254118 137748 254124 137760
rect 251324 137720 254124 137748
rect 251324 137708 251330 137720
rect 254118 137708 254124 137720
rect 254176 137708 254182 137760
rect 323578 137300 323584 137352
rect 323636 137340 323642 137352
rect 324406 137340 324412 137352
rect 323636 137312 324412 137340
rect 323636 137300 323642 137312
rect 324406 137300 324412 137312
rect 324464 137300 324470 137352
rect 187050 137232 187056 137284
rect 187108 137272 187114 137284
rect 214466 137272 214472 137284
rect 187108 137244 214472 137272
rect 187108 137232 187114 137244
rect 214466 137232 214472 137244
rect 214524 137232 214530 137284
rect 266998 136756 267004 136808
rect 267056 136796 267062 136808
rect 307478 136796 307484 136808
rect 267056 136768 307484 136796
rect 267056 136756 267062 136768
rect 307478 136756 307484 136768
rect 307536 136756 307542 136808
rect 250622 136688 250628 136740
rect 250680 136728 250686 136740
rect 307570 136728 307576 136740
rect 250680 136700 307576 136728
rect 250680 136688 250686 136700
rect 307570 136688 307576 136700
rect 307628 136688 307634 136740
rect 169110 136620 169116 136672
rect 169168 136660 169174 136672
rect 214098 136660 214104 136672
rect 169168 136632 214104 136660
rect 169168 136620 169174 136632
rect 214098 136620 214104 136632
rect 214156 136620 214162 136672
rect 250438 136620 250444 136672
rect 250496 136660 250502 136672
rect 307662 136660 307668 136672
rect 250496 136632 307668 136660
rect 250496 136620 250502 136632
rect 307662 136620 307668 136632
rect 307720 136620 307726 136672
rect 252462 136552 252468 136604
rect 252520 136592 252526 136604
rect 294598 136592 294604 136604
rect 252520 136564 294604 136592
rect 252520 136552 252526 136564
rect 294598 136552 294604 136564
rect 294656 136552 294662 136604
rect 252094 136484 252100 136536
rect 252152 136524 252158 136536
rect 265894 136524 265900 136536
rect 252152 136496 265900 136524
rect 252152 136484 252158 136496
rect 265894 136484 265900 136496
rect 265952 136484 265958 136536
rect 252186 135940 252192 135992
rect 252244 135980 252250 135992
rect 278130 135980 278136 135992
rect 252244 135952 278136 135980
rect 252244 135940 252250 135952
rect 278130 135940 278136 135952
rect 278188 135940 278194 135992
rect 264882 135872 264888 135924
rect 264940 135912 264946 135924
rect 302234 135912 302240 135924
rect 264940 135884 302240 135912
rect 264940 135872 264946 135884
rect 302234 135872 302240 135884
rect 302292 135872 302298 135924
rect 302878 135396 302884 135448
rect 302936 135436 302942 135448
rect 307478 135436 307484 135448
rect 302936 135408 307484 135436
rect 302936 135396 302942 135408
rect 307478 135396 307484 135408
rect 307536 135396 307542 135448
rect 172054 135328 172060 135380
rect 172112 135368 172118 135380
rect 214006 135368 214012 135380
rect 172112 135340 214012 135368
rect 172112 135328 172118 135340
rect 214006 135328 214012 135340
rect 214064 135328 214070 135380
rect 294690 135328 294696 135380
rect 294748 135368 294754 135380
rect 307662 135368 307668 135380
rect 294748 135340 307668 135368
rect 294748 135328 294754 135340
rect 307662 135328 307668 135340
rect 307720 135328 307726 135380
rect 169018 135260 169024 135312
rect 169076 135300 169082 135312
rect 213914 135300 213920 135312
rect 169076 135272 213920 135300
rect 169076 135260 169082 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 278314 135260 278320 135312
rect 278372 135300 278378 135312
rect 306926 135300 306932 135312
rect 278372 135272 306932 135300
rect 278372 135260 278378 135272
rect 306926 135260 306932 135272
rect 306984 135260 306990 135312
rect 252462 135192 252468 135244
rect 252520 135232 252526 135244
rect 283650 135232 283656 135244
rect 252520 135204 283656 135232
rect 252520 135192 252526 135204
rect 283650 135192 283656 135204
rect 283708 135192 283714 135244
rect 324314 135192 324320 135244
rect 324372 135232 324378 135244
rect 350626 135232 350632 135244
rect 324372 135204 350632 135232
rect 324372 135192 324378 135204
rect 350626 135192 350632 135204
rect 350684 135192 350690 135244
rect 252278 135124 252284 135176
rect 252336 135164 252342 135176
rect 269758 135164 269764 135176
rect 252336 135136 269764 135164
rect 252336 135124 252342 135136
rect 269758 135124 269764 135136
rect 269816 135124 269822 135176
rect 324498 135124 324504 135176
rect 324556 135164 324562 135176
rect 342438 135164 342444 135176
rect 324556 135136 342444 135164
rect 324556 135124 324562 135136
rect 342438 135124 342444 135136
rect 342496 135124 342502 135176
rect 269942 134512 269948 134564
rect 270000 134552 270006 134564
rect 307294 134552 307300 134564
rect 270000 134524 307300 134552
rect 270000 134512 270006 134524
rect 307294 134512 307300 134524
rect 307352 134512 307358 134564
rect 279510 134036 279516 134088
rect 279568 134076 279574 134088
rect 307478 134076 307484 134088
rect 279568 134048 307484 134076
rect 279568 134036 279574 134048
rect 307478 134036 307484 134048
rect 307536 134036 307542 134088
rect 295978 133968 295984 134020
rect 296036 134008 296042 134020
rect 307662 134008 307668 134020
rect 296036 133980 307668 134008
rect 296036 133968 296042 133980
rect 307662 133968 307668 133980
rect 307720 133968 307726 134020
rect 166258 133900 166264 133952
rect 166316 133940 166322 133952
rect 213914 133940 213920 133952
rect 166316 133912 213920 133940
rect 166316 133900 166322 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 251266 133832 251272 133884
rect 251324 133872 251330 133884
rect 281074 133872 281080 133884
rect 251324 133844 281080 133872
rect 251324 133832 251330 133844
rect 281074 133832 281080 133844
rect 281132 133832 281138 133884
rect 324314 133832 324320 133884
rect 324372 133872 324378 133884
rect 331306 133872 331312 133884
rect 324372 133844 331312 133872
rect 324372 133832 324378 133844
rect 331306 133832 331312 133844
rect 331364 133832 331370 133884
rect 252462 133764 252468 133816
rect 252520 133804 252526 133816
rect 265710 133804 265716 133816
rect 252520 133776 265716 133804
rect 252520 133764 252526 133776
rect 265710 133764 265716 133776
rect 265768 133764 265774 133816
rect 252370 133696 252376 133748
rect 252428 133736 252434 133748
rect 262950 133736 262956 133748
rect 252428 133708 262956 133736
rect 252428 133696 252434 133708
rect 262950 133696 262956 133708
rect 263008 133696 263014 133748
rect 280798 133220 280804 133272
rect 280856 133260 280862 133272
rect 298094 133260 298100 133272
rect 280856 133232 298100 133260
rect 280856 133220 280862 133232
rect 298094 133220 298100 133232
rect 298152 133220 298158 133272
rect 263134 133152 263140 133204
rect 263192 133192 263198 133204
rect 307110 133192 307116 133204
rect 263192 133164 307116 133192
rect 263192 133152 263198 133164
rect 307110 133152 307116 133164
rect 307168 133152 307174 133204
rect 301590 132608 301596 132660
rect 301648 132648 301654 132660
rect 307662 132648 307668 132660
rect 301648 132620 307668 132648
rect 301648 132608 301654 132620
rect 307662 132608 307668 132620
rect 307720 132608 307726 132660
rect 282270 132540 282276 132592
rect 282328 132580 282334 132592
rect 306926 132580 306932 132592
rect 282328 132552 306932 132580
rect 282328 132540 282334 132552
rect 306926 132540 306932 132552
rect 306984 132540 306990 132592
rect 173158 132472 173164 132524
rect 173216 132512 173222 132524
rect 213914 132512 213920 132524
rect 173216 132484 213920 132512
rect 173216 132472 173222 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 280982 132472 280988 132524
rect 281040 132512 281046 132524
rect 306558 132512 306564 132524
rect 281040 132484 306564 132512
rect 281040 132472 281046 132484
rect 306558 132472 306564 132484
rect 306616 132472 306622 132524
rect 251726 132404 251732 132456
rect 251784 132444 251790 132456
rect 304258 132444 304264 132456
rect 251784 132416 304264 132444
rect 251784 132404 251790 132416
rect 304258 132404 304264 132416
rect 304316 132404 304322 132456
rect 324314 132404 324320 132456
rect 324372 132444 324378 132456
rect 354766 132444 354772 132456
rect 324372 132416 354772 132444
rect 324372 132404 324378 132416
rect 354766 132404 354772 132416
rect 354824 132404 354830 132456
rect 252278 132336 252284 132388
rect 252336 132376 252342 132388
rect 258902 132376 258908 132388
rect 252336 132348 258908 132376
rect 252336 132336 252342 132348
rect 258902 132336 258908 132348
rect 258960 132336 258966 132388
rect 252002 131724 252008 131776
rect 252060 131764 252066 131776
rect 285122 131764 285128 131776
rect 252060 131736 285128 131764
rect 252060 131724 252066 131736
rect 285122 131724 285128 131736
rect 285180 131724 285186 131776
rect 285030 131180 285036 131232
rect 285088 131220 285094 131232
rect 307662 131220 307668 131232
rect 285088 131192 307668 131220
rect 285088 131180 285094 131192
rect 307662 131180 307668 131192
rect 307720 131180 307726 131232
rect 283834 131112 283840 131164
rect 283892 131152 283898 131164
rect 306926 131152 306932 131164
rect 283892 131124 306932 131152
rect 283892 131112 283898 131124
rect 306926 131112 306932 131124
rect 306984 131112 306990 131164
rect 252278 131044 252284 131096
rect 252336 131084 252342 131096
rect 279418 131084 279424 131096
rect 252336 131056 279424 131084
rect 252336 131044 252342 131056
rect 279418 131044 279424 131056
rect 279476 131044 279482 131096
rect 324314 131044 324320 131096
rect 324372 131084 324378 131096
rect 343818 131084 343824 131096
rect 324372 131056 343824 131084
rect 324372 131044 324378 131056
rect 343818 131044 343824 131056
rect 343876 131044 343882 131096
rect 252370 130976 252376 131028
rect 252428 131016 252434 131028
rect 273898 131016 273904 131028
rect 252428 130988 273904 131016
rect 252428 130976 252434 130988
rect 273898 130976 273904 130988
rect 273956 130976 273962 131028
rect 252462 130908 252468 130960
rect 252520 130948 252526 130960
rect 267182 130948 267188 130960
rect 252520 130920 267188 130948
rect 252520 130908 252526 130920
rect 267182 130908 267188 130920
rect 267240 130908 267246 130960
rect 256694 130364 256700 130416
rect 256752 130404 256758 130416
rect 305086 130404 305092 130416
rect 256752 130376 305092 130404
rect 256752 130364 256758 130376
rect 305086 130364 305092 130376
rect 305144 130364 305150 130416
rect 174538 129820 174544 129872
rect 174596 129860 174602 129872
rect 213914 129860 213920 129872
rect 174596 129832 213920 129860
rect 174596 129820 174602 129832
rect 213914 129820 213920 129832
rect 213972 129820 213978 129872
rect 278222 129820 278228 129872
rect 278280 129860 278286 129872
rect 307294 129860 307300 129872
rect 278280 129832 307300 129860
rect 278280 129820 278286 129832
rect 307294 129820 307300 129832
rect 307352 129820 307358 129872
rect 171870 129752 171876 129804
rect 171928 129792 171934 129804
rect 214006 129792 214012 129804
rect 171928 129764 214012 129792
rect 171928 129752 171934 129764
rect 214006 129752 214012 129764
rect 214064 129752 214070 129804
rect 273990 129752 273996 129804
rect 274048 129792 274054 129804
rect 307662 129792 307668 129804
rect 274048 129764 307668 129792
rect 274048 129752 274054 129764
rect 307662 129752 307668 129764
rect 307720 129752 307726 129804
rect 252462 129684 252468 129736
rect 252520 129724 252526 129736
rect 287882 129724 287888 129736
rect 252520 129696 287888 129724
rect 252520 129684 252526 129696
rect 287882 129684 287888 129696
rect 287940 129684 287946 129736
rect 324406 129684 324412 129736
rect 324464 129724 324470 129736
rect 329834 129724 329840 129736
rect 324464 129696 329840 129724
rect 324464 129684 324470 129696
rect 329834 129684 329840 129696
rect 329892 129684 329898 129736
rect 252370 129616 252376 129668
rect 252428 129656 252434 129668
rect 264330 129656 264336 129668
rect 252428 129628 264336 129656
rect 252428 129616 252434 129628
rect 264330 129616 264336 129628
rect 264388 129616 264394 129668
rect 324314 129616 324320 129668
rect 324372 129656 324378 129668
rect 330018 129656 330024 129668
rect 324372 129628 330024 129656
rect 324372 129616 324378 129628
rect 330018 129616 330024 129628
rect 330076 129616 330082 129668
rect 252278 129548 252284 129600
rect 252336 129588 252342 129600
rect 261478 129588 261484 129600
rect 252336 129560 261484 129588
rect 252336 129548 252342 129560
rect 261478 129548 261484 129560
rect 261536 129548 261542 129600
rect 287790 128460 287796 128512
rect 287848 128500 287854 128512
rect 307662 128500 307668 128512
rect 287848 128472 307668 128500
rect 287848 128460 287854 128472
rect 307662 128460 307668 128472
rect 307720 128460 307726 128512
rect 286318 128392 286324 128444
rect 286376 128432 286382 128444
rect 307294 128432 307300 128444
rect 286376 128404 307300 128432
rect 286376 128392 286382 128404
rect 307294 128392 307300 128404
rect 307352 128392 307358 128444
rect 188338 128324 188344 128376
rect 188396 128364 188402 128376
rect 213914 128364 213920 128376
rect 188396 128336 213920 128364
rect 188396 128324 188402 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 269850 128324 269856 128376
rect 269908 128364 269914 128376
rect 306742 128364 306748 128376
rect 269908 128336 306748 128364
rect 269908 128324 269914 128336
rect 306742 128324 306748 128336
rect 306800 128324 306806 128376
rect 251818 128256 251824 128308
rect 251876 128296 251882 128308
rect 282362 128296 282368 128308
rect 251876 128268 282368 128296
rect 251876 128256 251882 128268
rect 282362 128256 282368 128268
rect 282420 128256 282426 128308
rect 324406 128256 324412 128308
rect 324464 128296 324470 128308
rect 347958 128296 347964 128308
rect 324464 128268 347964 128296
rect 324464 128256 324470 128268
rect 347958 128256 347964 128268
rect 348016 128256 348022 128308
rect 252462 128188 252468 128240
rect 252520 128228 252526 128240
rect 267090 128228 267096 128240
rect 252520 128200 267096 128228
rect 252520 128188 252526 128200
rect 267090 128188 267096 128200
rect 267148 128188 267154 128240
rect 324314 128188 324320 128240
rect 324372 128228 324378 128240
rect 329926 128228 329932 128240
rect 324372 128200 329932 128228
rect 324372 128188 324378 128200
rect 329926 128188 329932 128200
rect 329984 128188 329990 128240
rect 252370 128120 252376 128172
rect 252428 128160 252434 128172
rect 263042 128160 263048 128172
rect 252428 128132 263048 128160
rect 252428 128120 252434 128132
rect 263042 128120 263048 128132
rect 263100 128120 263106 128172
rect 171778 127576 171784 127628
rect 171836 127616 171842 127628
rect 210602 127616 210608 127628
rect 171836 127588 210608 127616
rect 171836 127576 171842 127588
rect 210602 127576 210608 127588
rect 210660 127576 210666 127628
rect 294782 127576 294788 127628
rect 294840 127616 294846 127628
rect 307202 127616 307208 127628
rect 294840 127588 307208 127616
rect 294840 127576 294846 127588
rect 307202 127576 307208 127588
rect 307260 127576 307266 127628
rect 189810 127032 189816 127084
rect 189868 127072 189874 127084
rect 213914 127072 213920 127084
rect 189868 127044 213920 127072
rect 189868 127032 189874 127044
rect 213914 127032 213920 127044
rect 213972 127032 213978 127084
rect 279418 127032 279424 127084
rect 279476 127072 279482 127084
rect 307570 127072 307576 127084
rect 279476 127044 307576 127072
rect 279476 127032 279482 127044
rect 307570 127032 307576 127044
rect 307628 127032 307634 127084
rect 171962 126964 171968 127016
rect 172020 127004 172026 127016
rect 214006 127004 214012 127016
rect 172020 126976 214012 127004
rect 172020 126964 172026 126976
rect 214006 126964 214012 126976
rect 214064 126964 214070 127016
rect 271138 126964 271144 127016
rect 271196 127004 271202 127016
rect 307662 127004 307668 127016
rect 271196 126976 307668 127004
rect 271196 126964 271202 126976
rect 307662 126964 307668 126976
rect 307720 126964 307726 127016
rect 252186 126896 252192 126948
rect 252244 126936 252250 126948
rect 271230 126936 271236 126948
rect 252244 126908 271236 126936
rect 252244 126896 252250 126908
rect 271230 126896 271236 126908
rect 271288 126896 271294 126948
rect 324314 126896 324320 126948
rect 324372 126936 324378 126948
rect 342530 126936 342536 126948
rect 324372 126908 342536 126936
rect 324372 126896 324378 126908
rect 342530 126896 342536 126908
rect 342588 126896 342594 126948
rect 449158 126896 449164 126948
rect 449216 126936 449222 126948
rect 580166 126936 580172 126948
rect 449216 126908 580172 126936
rect 449216 126896 449222 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 252462 126692 252468 126744
rect 252520 126732 252526 126744
rect 257522 126732 257528 126744
rect 252520 126704 257528 126732
rect 252520 126692 252526 126704
rect 257522 126692 257528 126704
rect 257580 126692 257586 126744
rect 276014 126284 276020 126336
rect 276072 126324 276078 126336
rect 292022 126324 292028 126336
rect 276072 126296 292028 126324
rect 276072 126284 276078 126296
rect 292022 126284 292028 126296
rect 292080 126284 292086 126336
rect 251542 126216 251548 126268
rect 251600 126256 251606 126268
rect 305638 126256 305644 126268
rect 251600 126228 305644 126256
rect 251600 126216 251606 126228
rect 305638 126216 305644 126228
rect 305696 126216 305702 126268
rect 211982 125672 211988 125724
rect 212040 125712 212046 125724
rect 214742 125712 214748 125724
rect 212040 125684 214748 125712
rect 212040 125672 212046 125684
rect 214742 125672 214748 125684
rect 214800 125672 214806 125724
rect 289170 125672 289176 125724
rect 289228 125712 289234 125724
rect 306558 125712 306564 125724
rect 289228 125684 306564 125712
rect 289228 125672 289234 125684
rect 306558 125672 306564 125684
rect 306616 125672 306622 125724
rect 166350 125604 166356 125656
rect 166408 125644 166414 125656
rect 213914 125644 213920 125656
rect 166408 125616 213920 125644
rect 166408 125604 166414 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 260282 125604 260288 125656
rect 260340 125644 260346 125656
rect 306926 125644 306932 125656
rect 260340 125616 306932 125644
rect 260340 125604 260346 125616
rect 306926 125604 306932 125616
rect 306984 125604 306990 125656
rect 252462 125060 252468 125112
rect 252520 125100 252526 125112
rect 258994 125100 259000 125112
rect 252520 125072 259000 125100
rect 252520 125060 252526 125072
rect 258994 125060 259000 125072
rect 259052 125060 259058 125112
rect 252186 124856 252192 124908
rect 252244 124896 252250 124908
rect 301498 124896 301504 124908
rect 252244 124868 301504 124896
rect 252244 124856 252250 124868
rect 301498 124856 301504 124868
rect 301556 124856 301562 124908
rect 252462 124584 252468 124636
rect 252520 124624 252526 124636
rect 260190 124624 260196 124636
rect 252520 124596 260196 124624
rect 252520 124584 252526 124596
rect 260190 124584 260196 124596
rect 260248 124584 260254 124636
rect 264330 124380 264336 124432
rect 264388 124420 264394 124432
rect 306926 124420 306932 124432
rect 264388 124392 306932 124420
rect 264388 124380 264394 124392
rect 306926 124380 306932 124392
rect 306984 124380 306990 124432
rect 184382 124244 184388 124296
rect 184440 124284 184446 124296
rect 214006 124284 214012 124296
rect 184440 124256 214012 124284
rect 184440 124244 184446 124256
rect 214006 124244 214012 124256
rect 214064 124244 214070 124296
rect 265710 124244 265716 124296
rect 265768 124284 265774 124296
rect 307662 124284 307668 124296
rect 265768 124256 307668 124284
rect 265768 124244 265774 124256
rect 307662 124244 307668 124256
rect 307720 124244 307726 124296
rect 167730 124176 167736 124228
rect 167788 124216 167794 124228
rect 213914 124216 213920 124228
rect 167788 124188 213920 124216
rect 167788 124176 167794 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 301774 124176 301780 124228
rect 301832 124216 301838 124228
rect 307478 124216 307484 124228
rect 301832 124188 307484 124216
rect 301832 124176 301838 124188
rect 307478 124176 307484 124188
rect 307536 124176 307542 124228
rect 252462 124108 252468 124160
rect 252520 124148 252526 124160
rect 290642 124148 290648 124160
rect 252520 124120 290648 124148
rect 252520 124108 252526 124120
rect 290642 124108 290648 124120
rect 290700 124108 290706 124160
rect 324314 124108 324320 124160
rect 324372 124148 324378 124160
rect 334158 124148 334164 124160
rect 324372 124120 334164 124148
rect 324372 124108 324378 124120
rect 334158 124108 334164 124120
rect 334216 124108 334222 124160
rect 251266 124040 251272 124092
rect 251324 124080 251330 124092
rect 268470 124080 268476 124092
rect 251324 124052 268476 124080
rect 251324 124040 251330 124052
rect 268470 124040 268476 124052
rect 268528 124040 268534 124092
rect 251818 123428 251824 123480
rect 251876 123468 251882 123480
rect 284938 123468 284944 123480
rect 251876 123440 284944 123468
rect 251876 123428 251882 123440
rect 284938 123428 284944 123440
rect 284996 123428 285002 123480
rect 290458 122952 290464 123004
rect 290516 122992 290522 123004
rect 307570 122992 307576 123004
rect 290516 122964 307576 122992
rect 290516 122952 290522 122964
rect 307570 122952 307576 122964
rect 307628 122952 307634 123004
rect 176010 122884 176016 122936
rect 176068 122924 176074 122936
rect 214006 122924 214012 122936
rect 176068 122896 214012 122924
rect 176068 122884 176074 122896
rect 214006 122884 214012 122896
rect 214064 122884 214070 122936
rect 287882 122884 287888 122936
rect 287940 122924 287946 122936
rect 307662 122924 307668 122936
rect 287940 122896 307668 122924
rect 287940 122884 287946 122896
rect 307662 122884 307668 122896
rect 307720 122884 307726 122936
rect 170490 122816 170496 122868
rect 170548 122856 170554 122868
rect 213914 122856 213920 122868
rect 170548 122828 213920 122856
rect 170548 122816 170554 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 285122 122816 285128 122868
rect 285180 122856 285186 122868
rect 307478 122856 307484 122868
rect 285180 122828 307484 122856
rect 285180 122816 285186 122828
rect 307478 122816 307484 122828
rect 307536 122816 307542 122868
rect 252462 122748 252468 122800
rect 252520 122788 252526 122800
rect 298738 122788 298744 122800
rect 252520 122760 298744 122788
rect 252520 122748 252526 122760
rect 298738 122748 298744 122760
rect 298796 122748 298802 122800
rect 324314 122748 324320 122800
rect 324372 122788 324378 122800
rect 351914 122788 351920 122800
rect 324372 122760 351920 122788
rect 324372 122748 324378 122760
rect 351914 122748 351920 122760
rect 351972 122748 351978 122800
rect 252370 122680 252376 122732
rect 252428 122720 252434 122732
rect 261754 122720 261760 122732
rect 252428 122692 261760 122720
rect 252428 122680 252434 122692
rect 261754 122680 261760 122692
rect 261812 122680 261818 122732
rect 324406 122680 324412 122732
rect 324464 122720 324470 122732
rect 343726 122720 343732 122732
rect 324464 122692 343732 122720
rect 324464 122680 324470 122692
rect 343726 122680 343732 122692
rect 343784 122680 343790 122732
rect 251726 122612 251732 122664
rect 251784 122652 251790 122664
rect 258810 122652 258816 122664
rect 251784 122624 258816 122652
rect 251784 122612 251790 122624
rect 258810 122612 258816 122624
rect 258868 122612 258874 122664
rect 173342 122068 173348 122120
rect 173400 122108 173406 122120
rect 214742 122108 214748 122120
rect 173400 122080 214748 122108
rect 173400 122068 173406 122080
rect 214742 122068 214748 122080
rect 214800 122068 214806 122120
rect 300210 121592 300216 121644
rect 300268 121632 300274 121644
rect 307478 121632 307484 121644
rect 300268 121604 307484 121632
rect 300268 121592 300274 121604
rect 307478 121592 307484 121604
rect 307536 121592 307542 121644
rect 210510 121524 210516 121576
rect 210568 121564 210574 121576
rect 214006 121564 214012 121576
rect 210568 121536 214012 121564
rect 210568 121524 210574 121536
rect 214006 121524 214012 121536
rect 214064 121524 214070 121576
rect 283650 121524 283656 121576
rect 283708 121564 283714 121576
rect 307662 121564 307668 121576
rect 283708 121536 307668 121564
rect 283708 121524 283714 121536
rect 307662 121524 307668 121536
rect 307720 121524 307726 121576
rect 188430 121456 188436 121508
rect 188488 121496 188494 121508
rect 213914 121496 213920 121508
rect 188488 121468 213920 121496
rect 188488 121456 188494 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 261478 121456 261484 121508
rect 261536 121496 261542 121508
rect 306926 121496 306932 121508
rect 261536 121468 306932 121496
rect 261536 121456 261542 121468
rect 306926 121456 306932 121468
rect 306984 121456 306990 121508
rect 252370 121388 252376 121440
rect 252428 121428 252434 121440
rect 302970 121428 302976 121440
rect 252428 121400 302976 121428
rect 252428 121388 252434 121400
rect 302970 121388 302976 121400
rect 303028 121388 303034 121440
rect 324406 121388 324412 121440
rect 324464 121428 324470 121440
rect 339678 121428 339684 121440
rect 324464 121400 339684 121428
rect 324464 121388 324470 121400
rect 339678 121388 339684 121400
rect 339736 121388 339742 121440
rect 252462 121320 252468 121372
rect 252520 121360 252526 121372
rect 283742 121360 283748 121372
rect 252520 121332 283748 121360
rect 252520 121320 252526 121332
rect 283742 121320 283748 121332
rect 283800 121320 283806 121372
rect 251726 121252 251732 121304
rect 251784 121292 251790 121304
rect 260098 121292 260104 121304
rect 251784 121264 260104 121292
rect 251784 121252 251790 121264
rect 260098 121252 260104 121264
rect 260156 121252 260162 121304
rect 324314 120980 324320 121032
rect 324372 121020 324378 121032
rect 327074 121020 327080 121032
rect 324372 120992 327080 121020
rect 324372 120980 324378 120992
rect 327074 120980 327080 120992
rect 327132 120980 327138 121032
rect 171778 120708 171784 120760
rect 171836 120748 171842 120760
rect 214926 120748 214932 120760
rect 171836 120720 214932 120748
rect 171836 120708 171842 120720
rect 214926 120708 214932 120720
rect 214984 120708 214990 120760
rect 304534 120232 304540 120284
rect 304592 120272 304598 120284
rect 307478 120272 307484 120284
rect 304592 120244 307484 120272
rect 304592 120232 304598 120244
rect 307478 120232 307484 120244
rect 307536 120232 307542 120284
rect 298922 120164 298928 120216
rect 298980 120204 298986 120216
rect 306742 120204 306748 120216
rect 298980 120176 306748 120204
rect 298980 120164 298986 120176
rect 306742 120164 306748 120176
rect 306800 120164 306806 120216
rect 196802 120096 196808 120148
rect 196860 120136 196866 120148
rect 213914 120136 213920 120148
rect 196860 120108 213920 120136
rect 196860 120096 196866 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 273898 120096 273904 120148
rect 273956 120136 273962 120148
rect 307662 120136 307668 120148
rect 273956 120108 307668 120136
rect 273956 120096 273962 120108
rect 307662 120096 307668 120108
rect 307720 120096 307726 120148
rect 252278 120028 252284 120080
rect 252336 120068 252342 120080
rect 265802 120068 265808 120080
rect 252336 120040 265808 120068
rect 252336 120028 252342 120040
rect 265802 120028 265808 120040
rect 265860 120028 265866 120080
rect 324314 120028 324320 120080
rect 324372 120068 324378 120080
rect 340966 120068 340972 120080
rect 324372 120040 340972 120068
rect 324372 120028 324378 120040
rect 340966 120028 340972 120040
rect 341024 120028 341030 120080
rect 251450 119960 251456 120012
rect 251508 120000 251514 120012
rect 254762 120000 254768 120012
rect 251508 119972 254768 120000
rect 251508 119960 251514 119972
rect 254762 119960 254768 119972
rect 254820 119960 254826 120012
rect 252094 119824 252100 119876
rect 252152 119864 252158 119876
rect 260374 119864 260380 119876
rect 252152 119836 260380 119864
rect 252152 119824 252158 119836
rect 260374 119824 260380 119836
rect 260432 119824 260438 119876
rect 260098 119348 260104 119400
rect 260156 119388 260162 119400
rect 307018 119388 307024 119400
rect 260156 119360 307024 119388
rect 260156 119348 260162 119360
rect 307018 119348 307024 119360
rect 307076 119348 307082 119400
rect 182910 118804 182916 118856
rect 182968 118844 182974 118856
rect 213914 118844 213920 118856
rect 182968 118816 213920 118844
rect 182968 118804 182974 118816
rect 213914 118804 213920 118816
rect 213972 118804 213978 118856
rect 301498 118804 301504 118856
rect 301556 118844 301562 118856
rect 306558 118844 306564 118856
rect 301556 118816 306564 118844
rect 301556 118804 301562 118816
rect 306558 118804 306564 118816
rect 306616 118804 306622 118856
rect 177482 118736 177488 118788
rect 177540 118776 177546 118788
rect 214006 118776 214012 118788
rect 177540 118748 214012 118776
rect 177540 118736 177546 118748
rect 214006 118736 214012 118748
rect 214064 118736 214070 118788
rect 293218 118736 293224 118788
rect 293276 118776 293282 118788
rect 307662 118776 307668 118788
rect 293276 118748 307668 118776
rect 293276 118736 293282 118748
rect 307662 118736 307668 118748
rect 307720 118736 307726 118788
rect 166442 118668 166448 118720
rect 166500 118708 166506 118720
rect 214098 118708 214104 118720
rect 166500 118680 214104 118708
rect 166500 118668 166506 118680
rect 214098 118668 214104 118680
rect 214156 118668 214162 118720
rect 269758 118668 269764 118720
rect 269816 118708 269822 118720
rect 306926 118708 306932 118720
rect 269816 118680 306932 118708
rect 269816 118668 269822 118680
rect 306926 118668 306932 118680
rect 306984 118668 306990 118720
rect 251726 118600 251732 118652
rect 251784 118640 251790 118652
rect 296070 118640 296076 118652
rect 251784 118612 296076 118640
rect 251784 118600 251790 118612
rect 296070 118600 296076 118612
rect 296128 118600 296134 118652
rect 324406 118600 324412 118652
rect 324464 118640 324470 118652
rect 347866 118640 347872 118652
rect 324464 118612 347872 118640
rect 324464 118600 324470 118612
rect 347866 118600 347872 118612
rect 347924 118600 347930 118652
rect 252462 118532 252468 118584
rect 252520 118572 252526 118584
rect 264422 118572 264428 118584
rect 252520 118544 264428 118572
rect 252520 118532 252526 118544
rect 264422 118532 264428 118544
rect 264480 118532 264486 118584
rect 324314 118532 324320 118584
rect 324372 118572 324378 118584
rect 339586 118572 339592 118584
rect 324372 118544 339592 118572
rect 324372 118532 324378 118544
rect 339586 118532 339592 118544
rect 339644 118532 339650 118584
rect 264974 117920 264980 117972
rect 265032 117960 265038 117972
rect 293126 117960 293132 117972
rect 265032 117932 293132 117960
rect 265032 117920 265038 117932
rect 293126 117920 293132 117932
rect 293184 117920 293190 117972
rect 252278 117852 252284 117904
rect 252336 117892 252342 117904
rect 257430 117892 257436 117904
rect 252336 117864 257436 117892
rect 252336 117852 252342 117864
rect 257430 117852 257436 117864
rect 257488 117852 257494 117904
rect 302970 117444 302976 117496
rect 303028 117484 303034 117496
rect 307570 117484 307576 117496
rect 303028 117456 307576 117484
rect 303028 117444 303034 117456
rect 307570 117444 307576 117456
rect 307628 117444 307634 117496
rect 185762 117376 185768 117428
rect 185820 117416 185826 117428
rect 214006 117416 214012 117428
rect 185820 117388 214012 117416
rect 185820 117376 185826 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 297450 117376 297456 117428
rect 297508 117416 297514 117428
rect 307662 117416 307668 117428
rect 297508 117388 307668 117416
rect 297508 117376 297514 117388
rect 307662 117376 307668 117388
rect 307720 117376 307726 117428
rect 167822 117308 167828 117360
rect 167880 117348 167886 117360
rect 213914 117348 213920 117360
rect 167880 117320 213920 117348
rect 167880 117308 167886 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 292022 117308 292028 117360
rect 292080 117348 292086 117360
rect 306558 117348 306564 117360
rect 292080 117320 306564 117348
rect 292080 117308 292086 117320
rect 306558 117308 306564 117320
rect 306616 117308 306622 117360
rect 251266 117240 251272 117292
rect 251324 117280 251330 117292
rect 278406 117280 278412 117292
rect 251324 117252 278412 117280
rect 251324 117240 251330 117252
rect 278406 117240 278412 117252
rect 278464 117240 278470 117292
rect 252462 117172 252468 117224
rect 252520 117212 252526 117224
rect 261570 117212 261576 117224
rect 252520 117184 261576 117212
rect 252520 117172 252526 117184
rect 261570 117172 261576 117184
rect 261628 117172 261634 117224
rect 282362 116084 282368 116136
rect 282420 116124 282426 116136
rect 307662 116124 307668 116136
rect 282420 116096 307668 116124
rect 282420 116084 282426 116096
rect 307662 116084 307668 116096
rect 307720 116084 307726 116136
rect 169294 116016 169300 116068
rect 169352 116056 169358 116068
rect 214006 116056 214012 116068
rect 169352 116028 214012 116056
rect 169352 116016 169358 116028
rect 214006 116016 214012 116028
rect 214064 116016 214070 116068
rect 278130 116016 278136 116068
rect 278188 116056 278194 116068
rect 306742 116056 306748 116068
rect 278188 116028 306748 116056
rect 278188 116016 278194 116028
rect 306742 116016 306748 116028
rect 306800 116016 306806 116068
rect 169202 115948 169208 116000
rect 169260 115988 169266 116000
rect 213914 115988 213920 116000
rect 169260 115960 213920 115988
rect 169260 115948 169266 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 262950 115948 262956 116000
rect 263008 115988 263014 116000
rect 307570 115988 307576 116000
rect 263008 115960 307576 115988
rect 263008 115948 263014 115960
rect 307570 115948 307576 115960
rect 307628 115948 307634 116000
rect 251542 115880 251548 115932
rect 251600 115920 251606 115932
rect 282454 115920 282460 115932
rect 251600 115892 282460 115920
rect 251600 115880 251606 115892
rect 282454 115880 282460 115892
rect 282512 115880 282518 115932
rect 324406 115880 324412 115932
rect 324464 115920 324470 115932
rect 354674 115920 354680 115932
rect 324464 115892 354680 115920
rect 324464 115880 324470 115892
rect 354674 115880 354680 115892
rect 354732 115880 354738 115932
rect 324314 115812 324320 115864
rect 324372 115852 324378 115864
rect 336734 115852 336740 115864
rect 324372 115824 336740 115852
rect 324372 115812 324378 115824
rect 336734 115812 336740 115824
rect 336792 115812 336798 115864
rect 251174 115608 251180 115660
rect 251232 115648 251238 115660
rect 253474 115648 253480 115660
rect 251232 115620 253480 115648
rect 251232 115608 251238 115620
rect 253474 115608 253480 115620
rect 253532 115608 253538 115660
rect 304442 114656 304448 114708
rect 304500 114696 304506 114708
rect 306742 114696 306748 114708
rect 304500 114668 306748 114696
rect 304500 114656 304506 114668
rect 306742 114656 306748 114668
rect 306800 114656 306806 114708
rect 203610 114588 203616 114640
rect 203668 114628 203674 114640
rect 214006 114628 214012 114640
rect 203668 114600 214012 114628
rect 203668 114588 203674 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 297634 114588 297640 114640
rect 297692 114628 297698 114640
rect 307570 114628 307576 114640
rect 297692 114600 307576 114628
rect 297692 114588 297698 114600
rect 307570 114588 307576 114600
rect 307628 114588 307634 114640
rect 173250 114520 173256 114572
rect 173308 114560 173314 114572
rect 213914 114560 213920 114572
rect 173308 114532 213920 114560
rect 173308 114520 173314 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 268470 114520 268476 114572
rect 268528 114560 268534 114572
rect 307662 114560 307668 114572
rect 268528 114532 307668 114560
rect 268528 114520 268534 114532
rect 307662 114520 307668 114532
rect 307720 114520 307726 114572
rect 252462 114452 252468 114504
rect 252520 114492 252526 114504
rect 285214 114492 285220 114504
rect 252520 114464 285220 114492
rect 252520 114452 252526 114464
rect 285214 114452 285220 114464
rect 285272 114452 285278 114504
rect 324314 114452 324320 114504
rect 324372 114492 324378 114504
rect 346486 114492 346492 114504
rect 324372 114464 346492 114492
rect 324372 114452 324378 114464
rect 346486 114452 346492 114464
rect 346544 114452 346550 114504
rect 252370 114384 252376 114436
rect 252428 114424 252434 114436
rect 276750 114424 276756 114436
rect 252428 114396 276756 114424
rect 252428 114384 252434 114396
rect 276750 114384 276756 114396
rect 276808 114384 276814 114436
rect 324406 114384 324412 114436
rect 324464 114424 324470 114436
rect 343634 114424 343640 114436
rect 324464 114396 343640 114424
rect 324464 114384 324470 114396
rect 343634 114384 343640 114396
rect 343692 114384 343698 114436
rect 252462 114316 252468 114368
rect 252520 114356 252526 114368
rect 261662 114356 261668 114368
rect 252520 114328 261668 114356
rect 252520 114316 252526 114328
rect 261662 114316 261668 114328
rect 261720 114316 261726 114368
rect 170766 113772 170772 113824
rect 170824 113812 170830 113824
rect 199378 113812 199384 113824
rect 170824 113784 199384 113812
rect 170824 113772 170830 113784
rect 199378 113772 199384 113784
rect 199436 113772 199442 113824
rect 177390 113228 177396 113280
rect 177448 113268 177454 113280
rect 213914 113268 213920 113280
rect 177448 113240 213920 113268
rect 177448 113228 177454 113240
rect 213914 113228 213920 113240
rect 213972 113228 213978 113280
rect 294598 113228 294604 113280
rect 294656 113268 294662 113280
rect 307662 113268 307668 113280
rect 294656 113240 307668 113268
rect 294656 113228 294662 113240
rect 307662 113228 307668 113240
rect 307720 113228 307726 113280
rect 170582 113160 170588 113212
rect 170640 113200 170646 113212
rect 214006 113200 214012 113212
rect 170640 113172 214012 113200
rect 170640 113160 170646 113172
rect 214006 113160 214012 113172
rect 214064 113160 214070 113212
rect 284938 113160 284944 113212
rect 284996 113200 285002 113212
rect 307570 113200 307576 113212
rect 284996 113172 307576 113200
rect 284996 113160 285002 113172
rect 307570 113160 307576 113172
rect 307628 113160 307634 113212
rect 324314 113092 324320 113144
rect 324372 113132 324378 113144
rect 332686 113132 332692 113144
rect 324372 113104 332692 113132
rect 324372 113092 324378 113104
rect 332686 113092 332692 113104
rect 332744 113092 332750 113144
rect 467098 113092 467104 113144
rect 467156 113132 467162 113144
rect 579798 113132 579804 113144
rect 467156 113104 579804 113132
rect 467156 113092 467162 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 251726 112956 251732 113008
rect 251784 112996 251790 113008
rect 255958 112996 255964 113008
rect 251784 112968 255964 112996
rect 251784 112956 251790 112968
rect 255958 112956 255964 112968
rect 256016 112956 256022 113008
rect 252094 112616 252100 112668
rect 252152 112656 252158 112668
rect 256326 112656 256332 112668
rect 252152 112628 256332 112656
rect 252152 112616 252158 112628
rect 256326 112616 256332 112628
rect 256384 112616 256390 112668
rect 252370 112412 252376 112464
rect 252428 112452 252434 112464
rect 299014 112452 299020 112464
rect 252428 112424 299020 112452
rect 252428 112412 252434 112424
rect 299014 112412 299020 112424
rect 299072 112412 299078 112464
rect 300302 111936 300308 111988
rect 300360 111976 300366 111988
rect 307662 111976 307668 111988
rect 300360 111948 307668 111976
rect 300360 111936 300366 111948
rect 307662 111936 307668 111948
rect 307720 111936 307726 111988
rect 207750 111868 207756 111920
rect 207808 111908 207814 111920
rect 214006 111908 214012 111920
rect 207808 111880 214012 111908
rect 207808 111868 207814 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 298830 111868 298836 111920
rect 298888 111908 298894 111920
rect 307478 111908 307484 111920
rect 298888 111880 307484 111908
rect 298888 111868 298894 111880
rect 307478 111868 307484 111880
rect 307536 111868 307542 111920
rect 189902 111800 189908 111852
rect 189960 111840 189966 111852
rect 213914 111840 213920 111852
rect 189960 111812 213920 111840
rect 189960 111800 189966 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 256050 111800 256056 111852
rect 256108 111840 256114 111852
rect 307570 111840 307576 111852
rect 256108 111812 307576 111840
rect 256108 111800 256114 111812
rect 307570 111800 307576 111812
rect 307628 111800 307634 111852
rect 167914 111732 167920 111784
rect 167972 111772 167978 111784
rect 206370 111772 206376 111784
rect 167972 111744 206376 111772
rect 167972 111732 167978 111744
rect 206370 111732 206376 111744
rect 206428 111732 206434 111784
rect 252094 111732 252100 111784
rect 252152 111772 252158 111784
rect 275554 111772 275560 111784
rect 252152 111744 275560 111772
rect 252152 111732 252158 111744
rect 275554 111732 275560 111744
rect 275612 111732 275618 111784
rect 324314 111732 324320 111784
rect 324372 111772 324378 111784
rect 345014 111772 345020 111784
rect 324372 111744 345020 111772
rect 324372 111732 324378 111744
rect 345014 111732 345020 111744
rect 345072 111732 345078 111784
rect 324406 111664 324412 111716
rect 324464 111704 324470 111716
rect 334066 111704 334072 111716
rect 324464 111676 334072 111704
rect 324464 111664 324470 111676
rect 334066 111664 334072 111676
rect 334124 111664 334130 111716
rect 251634 111392 251640 111444
rect 251692 111432 251698 111444
rect 254670 111432 254676 111444
rect 251692 111404 254676 111432
rect 251692 111392 251698 111404
rect 254670 111392 254676 111404
rect 254728 111392 254734 111444
rect 251910 111052 251916 111104
rect 251968 111092 251974 111104
rect 279602 111092 279608 111104
rect 251968 111064 279608 111092
rect 251968 111052 251974 111064
rect 279602 111052 279608 111064
rect 279660 111052 279666 111104
rect 304258 110576 304264 110628
rect 304316 110616 304322 110628
rect 307662 110616 307668 110628
rect 304316 110588 307668 110616
rect 304316 110576 304322 110588
rect 307662 110576 307668 110588
rect 307720 110576 307726 110628
rect 200758 110508 200764 110560
rect 200816 110548 200822 110560
rect 214006 110548 214012 110560
rect 200816 110520 214012 110548
rect 200816 110508 200822 110520
rect 214006 110508 214012 110520
rect 214064 110508 214070 110560
rect 283742 110508 283748 110560
rect 283800 110548 283806 110560
rect 307478 110548 307484 110560
rect 283800 110520 307484 110548
rect 283800 110508 283806 110520
rect 307478 110508 307484 110520
rect 307536 110508 307542 110560
rect 184290 110440 184296 110492
rect 184348 110480 184354 110492
rect 213914 110480 213920 110492
rect 184348 110452 213920 110480
rect 184348 110440 184354 110452
rect 213914 110440 213920 110452
rect 213972 110440 213978 110492
rect 275370 110440 275376 110492
rect 275428 110480 275434 110492
rect 307570 110480 307576 110492
rect 275428 110452 307576 110480
rect 275428 110440 275434 110452
rect 307570 110440 307576 110452
rect 307628 110440 307634 110492
rect 168098 110372 168104 110424
rect 168156 110412 168162 110424
rect 177298 110412 177304 110424
rect 168156 110384 177304 110412
rect 168156 110372 168162 110384
rect 177298 110372 177304 110384
rect 177356 110372 177362 110424
rect 252094 110372 252100 110424
rect 252152 110412 252158 110424
rect 301682 110412 301688 110424
rect 252152 110384 301688 110412
rect 252152 110372 252158 110384
rect 301682 110372 301688 110384
rect 301740 110372 301746 110424
rect 324314 110372 324320 110424
rect 324372 110412 324378 110424
rect 339494 110412 339500 110424
rect 324372 110384 339500 110412
rect 324372 110372 324378 110384
rect 339494 110372 339500 110384
rect 339552 110372 339558 110424
rect 251542 110304 251548 110356
rect 251600 110344 251606 110356
rect 274174 110344 274180 110356
rect 251600 110316 274180 110344
rect 251600 110304 251606 110316
rect 274174 110304 274180 110316
rect 274232 110304 274238 110356
rect 252462 109488 252468 109540
rect 252520 109528 252526 109540
rect 258718 109528 258724 109540
rect 252520 109500 258724 109528
rect 252520 109488 252526 109500
rect 258718 109488 258724 109500
rect 258776 109488 258782 109540
rect 304350 109148 304356 109200
rect 304408 109188 304414 109200
rect 307478 109188 307484 109200
rect 304408 109160 307484 109188
rect 304408 109148 304414 109160
rect 307478 109148 307484 109160
rect 307536 109148 307542 109200
rect 178678 109080 178684 109132
rect 178736 109120 178742 109132
rect 214006 109120 214012 109132
rect 178736 109092 214012 109120
rect 178736 109080 178742 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 299014 109080 299020 109132
rect 299072 109120 299078 109132
rect 307570 109120 307576 109132
rect 299072 109092 307576 109120
rect 299072 109080 299078 109092
rect 307570 109080 307576 109092
rect 307628 109080 307634 109132
rect 168006 109012 168012 109064
rect 168064 109052 168070 109064
rect 213914 109052 213920 109064
rect 168064 109024 213920 109052
rect 168064 109012 168070 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 271230 109012 271236 109064
rect 271288 109052 271294 109064
rect 307662 109052 307668 109064
rect 271288 109024 307668 109052
rect 271288 109012 271294 109024
rect 307662 109012 307668 109024
rect 307720 109012 307726 109064
rect 167914 108944 167920 108996
rect 167972 108984 167978 108996
rect 184474 108984 184480 108996
rect 167972 108956 184480 108984
rect 167972 108944 167978 108956
rect 184474 108944 184480 108956
rect 184532 108944 184538 108996
rect 252002 108944 252008 108996
rect 252060 108984 252066 108996
rect 303154 108984 303160 108996
rect 252060 108956 303160 108984
rect 252060 108944 252066 108956
rect 303154 108944 303160 108956
rect 303212 108944 303218 108996
rect 252462 108876 252468 108928
rect 252520 108916 252526 108928
rect 276658 108916 276664 108928
rect 252520 108888 276664 108916
rect 252520 108876 252526 108888
rect 276658 108876 276664 108888
rect 276716 108876 276722 108928
rect 267090 107856 267096 107908
rect 267148 107896 267154 107908
rect 307662 107896 307668 107908
rect 267148 107868 307668 107896
rect 267148 107856 267154 107868
rect 307662 107856 307668 107868
rect 307720 107856 307726 107908
rect 205082 107720 205088 107772
rect 205140 107760 205146 107772
rect 213914 107760 213920 107772
rect 205140 107732 213920 107760
rect 205140 107720 205146 107732
rect 213914 107720 213920 107732
rect 213972 107720 213978 107772
rect 300394 107720 300400 107772
rect 300452 107760 300458 107772
rect 307570 107760 307576 107772
rect 300452 107732 307576 107760
rect 300452 107720 300458 107732
rect 307570 107720 307576 107732
rect 307628 107720 307634 107772
rect 188522 107652 188528 107704
rect 188580 107692 188586 107704
rect 214006 107692 214012 107704
rect 188580 107664 214012 107692
rect 188580 107652 188586 107664
rect 214006 107652 214012 107664
rect 214064 107652 214070 107704
rect 303062 107652 303068 107704
rect 303120 107692 303126 107704
rect 306926 107692 306932 107704
rect 303120 107664 306932 107692
rect 303120 107652 303126 107664
rect 306926 107652 306932 107664
rect 306984 107652 306990 107704
rect 251818 107584 251824 107636
rect 251876 107624 251882 107636
rect 272610 107624 272616 107636
rect 251876 107596 272616 107624
rect 251876 107584 251882 107596
rect 272610 107584 272616 107596
rect 272668 107584 272674 107636
rect 252094 107516 252100 107568
rect 252152 107556 252158 107568
rect 263134 107556 263140 107568
rect 252152 107528 263140 107556
rect 252152 107516 252158 107528
rect 263134 107516 263140 107528
rect 263192 107516 263198 107568
rect 252462 107448 252468 107500
rect 252520 107488 252526 107500
rect 257338 107488 257344 107500
rect 252520 107460 257344 107488
rect 252520 107448 252526 107460
rect 257338 107448 257344 107460
rect 257396 107448 257402 107500
rect 301682 106428 301688 106480
rect 301740 106468 301746 106480
rect 307478 106468 307484 106480
rect 301740 106440 307484 106468
rect 301740 106428 301746 106440
rect 307478 106428 307484 106440
rect 307536 106428 307542 106480
rect 192754 106360 192760 106412
rect 192812 106400 192818 106412
rect 213914 106400 213920 106412
rect 192812 106372 213920 106400
rect 192812 106360 192818 106372
rect 213914 106360 213920 106372
rect 213972 106360 213978 106412
rect 276658 106360 276664 106412
rect 276716 106400 276722 106412
rect 307570 106400 307576 106412
rect 276716 106372 307576 106400
rect 276716 106360 276722 106372
rect 307570 106360 307576 106372
rect 307628 106360 307634 106412
rect 174630 106292 174636 106344
rect 174688 106332 174694 106344
rect 214006 106332 214012 106344
rect 174688 106304 214012 106332
rect 174688 106292 174694 106304
rect 214006 106292 214012 106304
rect 214064 106292 214070 106344
rect 261570 106292 261576 106344
rect 261628 106332 261634 106344
rect 307662 106332 307668 106344
rect 261628 106304 307668 106332
rect 261628 106292 261634 106304
rect 307662 106292 307668 106304
rect 307720 106292 307726 106344
rect 252002 106224 252008 106276
rect 252060 106264 252066 106276
rect 299106 106264 299112 106276
rect 252060 106236 299112 106264
rect 252060 106224 252066 106236
rect 299106 106224 299112 106236
rect 299164 106224 299170 106276
rect 252278 106088 252284 106140
rect 252336 106128 252342 106140
rect 254578 106128 254584 106140
rect 252336 106100 254584 106128
rect 252336 106088 252342 106100
rect 254578 106088 254584 106100
rect 254636 106088 254642 106140
rect 252462 105748 252468 105800
rect 252520 105788 252526 105800
rect 256234 105788 256240 105800
rect 252520 105760 256240 105788
rect 252520 105748 252526 105760
rect 256234 105748 256240 105760
rect 256292 105748 256298 105800
rect 255958 105544 255964 105596
rect 256016 105584 256022 105596
rect 295334 105584 295340 105596
rect 256016 105556 295340 105584
rect 256016 105544 256022 105556
rect 295334 105544 295340 105556
rect 295392 105544 295398 105596
rect 212074 105000 212080 105052
rect 212132 105040 212138 105052
rect 214098 105040 214104 105052
rect 212132 105012 214104 105040
rect 212132 105000 212138 105012
rect 214098 105000 214104 105012
rect 214156 105000 214162 105052
rect 296070 105000 296076 105052
rect 296128 105040 296134 105052
rect 307478 105040 307484 105052
rect 296128 105012 307484 105040
rect 296128 105000 296134 105012
rect 307478 105000 307484 105012
rect 307536 105000 307542 105052
rect 206462 104932 206468 104984
rect 206520 104972 206526 104984
rect 213914 104972 213920 104984
rect 206520 104944 213920 104972
rect 206520 104932 206526 104944
rect 213914 104932 213920 104944
rect 213972 104932 213978 104984
rect 298738 104932 298744 104984
rect 298796 104972 298802 104984
rect 307662 104972 307668 104984
rect 298796 104944 307668 104972
rect 298796 104932 298802 104944
rect 307662 104932 307668 104944
rect 307720 104932 307726 104984
rect 194042 104864 194048 104916
rect 194100 104904 194106 104916
rect 214006 104904 214012 104916
rect 194100 104876 214012 104904
rect 194100 104864 194106 104876
rect 214006 104864 214012 104876
rect 214064 104864 214070 104916
rect 252462 104796 252468 104848
rect 252520 104836 252526 104848
rect 294782 104836 294788 104848
rect 252520 104808 294788 104836
rect 252520 104796 252526 104808
rect 294782 104796 294788 104808
rect 294840 104796 294846 104848
rect 324314 104796 324320 104848
rect 324372 104836 324378 104848
rect 328454 104836 328460 104848
rect 324372 104808 328460 104836
rect 324372 104796 324378 104808
rect 328454 104796 328460 104808
rect 328512 104796 328518 104848
rect 252186 104660 252192 104712
rect 252244 104700 252250 104712
rect 256142 104700 256148 104712
rect 252244 104672 256148 104700
rect 252244 104660 252250 104672
rect 256142 104660 256148 104672
rect 256200 104660 256206 104712
rect 251358 104116 251364 104168
rect 251416 104156 251422 104168
rect 287974 104156 287980 104168
rect 251416 104128 287980 104156
rect 251416 104116 251422 104128
rect 287974 104116 287980 104128
rect 288032 104116 288038 104168
rect 303154 103640 303160 103692
rect 303212 103680 303218 103692
rect 307570 103680 307576 103692
rect 303212 103652 307576 103680
rect 303212 103640 303218 103652
rect 307570 103640 307576 103652
rect 307628 103640 307634 103692
rect 206370 103572 206376 103624
rect 206428 103612 206434 103624
rect 214006 103612 214012 103624
rect 206428 103584 214012 103612
rect 206428 103572 206434 103584
rect 214006 103572 214012 103584
rect 214064 103572 214070 103624
rect 294874 103572 294880 103624
rect 294932 103612 294938 103624
rect 307662 103612 307668 103624
rect 294932 103584 307668 103612
rect 294932 103572 294938 103584
rect 307662 103572 307668 103584
rect 307720 103572 307726 103624
rect 177298 103504 177304 103556
rect 177356 103544 177362 103556
rect 213914 103544 213920 103556
rect 177356 103516 213920 103544
rect 177356 103504 177362 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 293310 103504 293316 103556
rect 293368 103544 293374 103556
rect 307478 103544 307484 103556
rect 293368 103516 307484 103544
rect 293368 103504 293374 103516
rect 307478 103504 307484 103516
rect 307536 103504 307542 103556
rect 252462 103436 252468 103488
rect 252520 103476 252526 103488
rect 262858 103476 262864 103488
rect 252520 103448 262864 103476
rect 252520 103436 252526 103448
rect 262858 103436 262864 103448
rect 262916 103436 262922 103488
rect 324314 103300 324320 103352
rect 324372 103340 324378 103352
rect 327258 103340 327264 103352
rect 324372 103312 327264 103340
rect 324372 103300 324378 103312
rect 327258 103300 327264 103312
rect 327316 103300 327322 103352
rect 170950 102756 170956 102808
rect 171008 102796 171014 102808
rect 204898 102796 204904 102808
rect 171008 102768 204904 102796
rect 171008 102756 171014 102768
rect 204898 102756 204904 102768
rect 204956 102756 204962 102808
rect 251174 102756 251180 102808
rect 251232 102796 251238 102808
rect 253382 102796 253388 102808
rect 251232 102768 253388 102796
rect 251232 102756 251238 102768
rect 253382 102756 253388 102768
rect 253440 102756 253446 102808
rect 293954 102796 293960 102808
rect 258046 102768 293960 102796
rect 251266 102688 251272 102740
rect 251324 102728 251330 102740
rect 258046 102728 258074 102768
rect 293954 102756 293960 102768
rect 294012 102756 294018 102808
rect 251324 102700 258074 102728
rect 251324 102688 251330 102700
rect 296162 102280 296168 102332
rect 296220 102320 296226 102332
rect 306742 102320 306748 102332
rect 296220 102292 306748 102320
rect 296220 102280 296226 102292
rect 306742 102280 306748 102292
rect 306800 102280 306806 102332
rect 294782 102212 294788 102264
rect 294840 102252 294846 102264
rect 307662 102252 307668 102264
rect 294840 102224 307668 102252
rect 294840 102212 294846 102224
rect 307662 102212 307668 102224
rect 307720 102212 307726 102264
rect 209222 102144 209228 102196
rect 209280 102184 209286 102196
rect 213914 102184 213920 102196
rect 209280 102156 213920 102184
rect 209280 102144 209286 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 261662 102144 261668 102196
rect 261720 102184 261726 102196
rect 307478 102184 307484 102196
rect 261720 102156 307484 102184
rect 261720 102144 261726 102156
rect 307478 102144 307484 102156
rect 307536 102144 307542 102196
rect 252462 102076 252468 102128
rect 252520 102116 252526 102128
rect 271322 102116 271328 102128
rect 252520 102088 271328 102116
rect 252520 102076 252526 102088
rect 271322 102076 271328 102088
rect 271380 102076 271386 102128
rect 324314 102076 324320 102128
rect 324372 102116 324378 102128
rect 349246 102116 349252 102128
rect 324372 102088 349252 102116
rect 324372 102076 324378 102088
rect 349246 102076 349252 102088
rect 349304 102076 349310 102128
rect 251174 101940 251180 101992
rect 251232 101980 251238 101992
rect 253290 101980 253296 101992
rect 251232 101952 253296 101980
rect 251232 101940 251238 101952
rect 253290 101940 253296 101952
rect 253348 101940 253354 101992
rect 170674 101396 170680 101448
rect 170732 101436 170738 101448
rect 214650 101436 214656 101448
rect 170732 101408 214656 101436
rect 170732 101396 170738 101408
rect 214650 101396 214656 101408
rect 214708 101396 214714 101448
rect 252186 101396 252192 101448
rect 252244 101436 252250 101448
rect 289078 101436 289084 101448
rect 252244 101408 289084 101436
rect 252244 101396 252250 101408
rect 289078 101396 289084 101408
rect 289136 101396 289142 101448
rect 292114 100784 292120 100836
rect 292172 100824 292178 100836
rect 306558 100824 306564 100836
rect 292172 100796 306564 100824
rect 292172 100784 292178 100796
rect 306558 100784 306564 100796
rect 306616 100784 306622 100836
rect 173434 100716 173440 100768
rect 173492 100756 173498 100768
rect 213914 100756 213920 100768
rect 173492 100728 213920 100756
rect 173492 100716 173498 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 250530 100716 250536 100768
rect 250588 100756 250594 100768
rect 307662 100756 307668 100768
rect 250588 100728 307668 100756
rect 250588 100716 250594 100728
rect 307662 100716 307668 100728
rect 307720 100716 307726 100768
rect 252002 100648 252008 100700
rect 252060 100688 252066 100700
rect 289354 100688 289360 100700
rect 252060 100660 289360 100688
rect 252060 100648 252066 100660
rect 289354 100648 289360 100660
rect 289412 100648 289418 100700
rect 512638 100648 512644 100700
rect 512696 100688 512702 100700
rect 580166 100688 580172 100700
rect 512696 100660 580172 100688
rect 512696 100648 512702 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 252462 100580 252468 100632
rect 252520 100620 252526 100632
rect 275462 100620 275468 100632
rect 252520 100592 275468 100620
rect 252520 100580 252526 100592
rect 275462 100580 275468 100592
rect 275520 100580 275526 100632
rect 251542 100512 251548 100564
rect 251600 100552 251606 100564
rect 269942 100552 269948 100564
rect 251600 100524 269948 100552
rect 251600 100512 251606 100524
rect 269942 100512 269948 100524
rect 270000 100512 270006 100564
rect 209130 99424 209136 99476
rect 209188 99464 209194 99476
rect 214006 99464 214012 99476
rect 209188 99436 214012 99464
rect 209188 99424 209194 99436
rect 214006 99424 214012 99436
rect 214064 99424 214070 99476
rect 289262 99424 289268 99476
rect 289320 99464 289326 99476
rect 307570 99464 307576 99476
rect 289320 99436 307576 99464
rect 289320 99424 289326 99436
rect 307570 99424 307576 99436
rect 307628 99424 307634 99476
rect 164878 99356 164884 99408
rect 164936 99396 164942 99408
rect 213914 99396 213920 99408
rect 164936 99368 213920 99396
rect 164936 99356 164942 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 274174 99356 274180 99408
rect 274232 99396 274238 99408
rect 307662 99396 307668 99408
rect 274232 99368 307668 99396
rect 274232 99356 274238 99368
rect 307662 99356 307668 99368
rect 307720 99356 307726 99408
rect 252462 98812 252468 98864
rect 252520 98852 252526 98864
rect 260098 98852 260104 98864
rect 252520 98824 260104 98852
rect 252520 98812 252526 98824
rect 260098 98812 260104 98824
rect 260156 98812 260162 98864
rect 293402 98132 293408 98184
rect 293460 98172 293466 98184
rect 307662 98172 307668 98184
rect 293460 98144 307668 98172
rect 293460 98132 293466 98144
rect 307662 98132 307668 98144
rect 307720 98132 307726 98184
rect 187142 98064 187148 98116
rect 187200 98104 187206 98116
rect 213914 98104 213920 98116
rect 187200 98076 213920 98104
rect 187200 98064 187206 98076
rect 213914 98064 213920 98076
rect 213972 98064 213978 98116
rect 260190 98064 260196 98116
rect 260248 98104 260254 98116
rect 307478 98104 307484 98116
rect 260248 98076 307484 98104
rect 260248 98064 260254 98076
rect 307478 98064 307484 98076
rect 307536 98064 307542 98116
rect 166534 97996 166540 98048
rect 166592 98036 166598 98048
rect 214006 98036 214012 98048
rect 166592 98008 214012 98036
rect 166592 97996 166598 98008
rect 214006 97996 214012 98008
rect 214064 97996 214070 98048
rect 256142 97996 256148 98048
rect 256200 98036 256206 98048
rect 307570 98036 307576 98048
rect 256200 98008 307576 98036
rect 256200 97996 256206 98008
rect 307570 97996 307576 98008
rect 307628 97996 307634 98048
rect 251174 97928 251180 97980
rect 251232 97968 251238 97980
rect 253198 97968 253204 97980
rect 251232 97940 253204 97968
rect 251232 97928 251238 97940
rect 253198 97928 253204 97940
rect 253256 97928 253262 97980
rect 289078 96772 289084 96824
rect 289136 96812 289142 96824
rect 306742 96812 306748 96824
rect 289136 96784 306748 96812
rect 289136 96772 289142 96784
rect 306742 96772 306748 96784
rect 306800 96772 306806 96824
rect 262858 96704 262864 96756
rect 262916 96744 262922 96756
rect 307662 96744 307668 96756
rect 262916 96716 307668 96744
rect 262916 96704 262922 96716
rect 307662 96704 307668 96716
rect 307720 96704 307726 96756
rect 193950 96636 193956 96688
rect 194008 96676 194014 96688
rect 213914 96676 213920 96688
rect 194008 96648 213920 96676
rect 194008 96636 194014 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 253290 96636 253296 96688
rect 253348 96676 253354 96688
rect 307478 96676 307484 96688
rect 253348 96648 307484 96676
rect 253348 96636 253354 96648
rect 307478 96636 307484 96648
rect 307536 96636 307542 96688
rect 258074 95888 258080 95940
rect 258132 95928 258138 95940
rect 283558 95928 283564 95940
rect 258132 95900 283564 95928
rect 258132 95888 258138 95900
rect 283558 95888 283564 95900
rect 283616 95888 283622 95940
rect 318058 95752 318064 95804
rect 318116 95792 318122 95804
rect 321462 95792 321468 95804
rect 318116 95764 321468 95792
rect 318116 95752 318122 95764
rect 321462 95752 321468 95764
rect 321520 95752 321526 95804
rect 185578 95140 185584 95192
rect 185636 95180 185642 95192
rect 323118 95180 323124 95192
rect 185636 95152 323124 95180
rect 185636 95140 185642 95152
rect 323118 95140 323124 95152
rect 323176 95140 323182 95192
rect 186958 95072 186964 95124
rect 187016 95112 187022 95124
rect 321646 95112 321652 95124
rect 187016 95084 321652 95112
rect 187016 95072 187022 95084
rect 321646 95072 321652 95084
rect 321704 95072 321710 95124
rect 199378 95004 199384 95056
rect 199436 95044 199442 95056
rect 321738 95044 321744 95056
rect 199436 95016 321744 95044
rect 199436 95004 199442 95016
rect 321738 95004 321744 95016
rect 321796 95004 321802 95056
rect 131942 94120 131948 94172
rect 132000 94160 132006 94172
rect 170398 94160 170404 94172
rect 132000 94132 170404 94160
rect 132000 94120 132006 94132
rect 170398 94120 170404 94132
rect 170456 94120 170462 94172
rect 151906 94052 151912 94104
rect 151964 94092 151970 94104
rect 195238 94092 195244 94104
rect 151964 94064 195244 94092
rect 151964 94052 151970 94064
rect 195238 94052 195244 94064
rect 195296 94052 195302 94104
rect 151722 93984 151728 94036
rect 151780 94024 151786 94036
rect 204990 94024 204996 94036
rect 151780 93996 204996 94024
rect 151780 93984 151786 93996
rect 204990 93984 204996 93996
rect 205048 93984 205054 94036
rect 109034 93916 109040 93968
rect 109092 93956 109098 93968
rect 169294 93956 169300 93968
rect 109092 93928 169300 93956
rect 109092 93916 109098 93928
rect 169294 93916 169300 93928
rect 169352 93916 169358 93968
rect 113726 93848 113732 93900
rect 113784 93888 113790 93900
rect 177482 93888 177488 93900
rect 113784 93860 177488 93888
rect 113784 93848 113790 93860
rect 177482 93848 177488 93860
rect 177540 93848 177546 93900
rect 241514 93848 241520 93900
rect 241572 93888 241578 93900
rect 250714 93888 250720 93900
rect 241572 93860 250720 93888
rect 241572 93848 241578 93860
rect 250714 93848 250720 93860
rect 250772 93848 250778 93900
rect 175918 93780 175924 93832
rect 175976 93820 175982 93832
rect 324498 93820 324504 93832
rect 175976 93792 324504 93820
rect 175976 93780 175982 93792
rect 324498 93780 324504 93792
rect 324556 93780 324562 93832
rect 63310 93712 63316 93764
rect 63368 93752 63374 93764
rect 209222 93752 209228 93764
rect 63368 93724 209228 93752
rect 63368 93712 63374 93724
rect 209222 93712 209228 93724
rect 209280 93712 209286 93764
rect 210602 93712 210608 93764
rect 210660 93752 210666 93764
rect 321554 93752 321560 93764
rect 210660 93724 321560 93752
rect 210660 93712 210666 93724
rect 321554 93712 321560 93724
rect 321612 93712 321618 93764
rect 64782 93644 64788 93696
rect 64840 93684 64846 93696
rect 206462 93684 206468 93696
rect 64840 93656 206468 93684
rect 64840 93644 64846 93656
rect 206462 93644 206468 93656
rect 206520 93644 206526 93696
rect 121730 93304 121736 93356
rect 121788 93344 121794 93356
rect 176010 93344 176016 93356
rect 121788 93316 176016 93344
rect 121788 93304 121794 93316
rect 176010 93304 176016 93316
rect 176068 93304 176074 93356
rect 124490 93236 124496 93288
rect 124548 93276 124554 93288
rect 182818 93276 182824 93288
rect 124548 93248 182824 93276
rect 124548 93236 124554 93248
rect 182818 93236 182824 93248
rect 182876 93236 182882 93288
rect 107746 93168 107752 93220
rect 107804 93208 107810 93220
rect 169202 93208 169208 93220
rect 107804 93180 169208 93208
rect 107804 93168 107810 93180
rect 169202 93168 169208 93180
rect 169260 93168 169266 93220
rect 102042 93100 102048 93152
rect 102100 93140 102106 93152
rect 174538 93140 174544 93152
rect 102100 93112 174544 93140
rect 102100 93100 102106 93112
rect 174538 93100 174544 93112
rect 174596 93100 174602 93152
rect 119338 92420 119344 92472
rect 119396 92460 119402 92472
rect 207658 92460 207664 92472
rect 119396 92432 207664 92460
rect 119396 92420 119402 92432
rect 207658 92420 207664 92432
rect 207716 92420 207722 92472
rect 120350 92352 120356 92404
rect 120408 92392 120414 92404
rect 181438 92392 181444 92404
rect 120408 92364 181444 92392
rect 120408 92352 120414 92364
rect 181438 92352 181444 92364
rect 181496 92352 181502 92404
rect 115474 92284 115480 92336
rect 115532 92324 115538 92336
rect 170674 92324 170680 92336
rect 115532 92296 170680 92324
rect 115532 92284 115538 92296
rect 170674 92284 170680 92296
rect 170732 92284 170738 92336
rect 133138 92216 133144 92268
rect 133196 92256 133202 92268
rect 187050 92256 187056 92268
rect 133196 92228 187056 92256
rect 133196 92216 133202 92228
rect 187050 92216 187056 92228
rect 187108 92216 187114 92268
rect 151722 92148 151728 92200
rect 151780 92188 151786 92200
rect 202138 92188 202144 92200
rect 151780 92160 202144 92188
rect 151780 92148 151786 92160
rect 202138 92148 202144 92160
rect 202196 92148 202202 92200
rect 125962 92080 125968 92132
rect 126020 92120 126026 92132
rect 171778 92120 171784 92132
rect 126020 92092 171784 92120
rect 126020 92080 126026 92092
rect 171778 92080 171784 92092
rect 171836 92080 171842 92132
rect 228358 91876 228364 91928
rect 228416 91916 228422 91928
rect 260282 91916 260288 91928
rect 228416 91888 260288 91916
rect 228416 91876 228422 91888
rect 260282 91876 260288 91888
rect 260340 91876 260346 91928
rect 192570 91808 192576 91860
rect 192628 91848 192634 91860
rect 232498 91848 232504 91860
rect 192628 91820 232504 91848
rect 192628 91808 192634 91820
rect 232498 91808 232504 91820
rect 232556 91808 232562 91860
rect 179138 91740 179144 91792
rect 179196 91780 179202 91792
rect 245654 91780 245660 91792
rect 179196 91752 245660 91780
rect 179196 91740 179202 91752
rect 245654 91740 245660 91752
rect 245712 91740 245718 91792
rect 94222 91264 94228 91316
rect 94280 91304 94286 91316
rect 120718 91304 120724 91316
rect 94280 91276 120724 91304
rect 94280 91264 94286 91276
rect 120718 91264 120724 91276
rect 120776 91264 120782 91316
rect 101858 91196 101864 91248
rect 101916 91236 101922 91248
rect 127618 91236 127624 91248
rect 101916 91208 127624 91236
rect 101916 91196 101922 91208
rect 127618 91196 127624 91208
rect 127676 91196 127682 91248
rect 85942 91128 85948 91180
rect 86000 91168 86006 91180
rect 120810 91168 120816 91180
rect 86000 91140 120816 91168
rect 86000 91128 86006 91140
rect 120810 91128 120816 91140
rect 120868 91128 120874 91180
rect 74810 91060 74816 91112
rect 74868 91100 74874 91112
rect 112438 91100 112444 91112
rect 74868 91072 112444 91100
rect 74868 91060 74874 91072
rect 112438 91060 112444 91072
rect 112496 91060 112502 91112
rect 67358 90992 67364 91044
rect 67416 91032 67422 91044
rect 214926 91032 214932 91044
rect 67416 91004 214932 91032
rect 67416 90992 67422 91004
rect 214926 90992 214932 91004
rect 214984 90992 214990 91044
rect 66162 90924 66168 90976
rect 66220 90964 66226 90976
rect 177298 90964 177304 90976
rect 66220 90936 177304 90964
rect 66220 90924 66226 90936
rect 177298 90924 177304 90936
rect 177356 90924 177362 90976
rect 196710 90924 196716 90976
rect 196768 90964 196774 90976
rect 323026 90964 323032 90976
rect 196768 90936 323032 90964
rect 196768 90924 196774 90936
rect 323026 90924 323032 90936
rect 323084 90924 323090 90976
rect 124122 90856 124128 90908
rect 124180 90896 124186 90908
rect 184382 90896 184388 90908
rect 124180 90868 184388 90896
rect 124180 90856 124186 90868
rect 184382 90856 184388 90868
rect 184440 90856 184446 90908
rect 115198 90788 115204 90840
rect 115256 90828 115262 90840
rect 166442 90828 166448 90840
rect 115256 90800 166448 90828
rect 115256 90788 115262 90800
rect 166442 90788 166448 90800
rect 166500 90788 166506 90840
rect 122834 90720 122840 90772
rect 122892 90760 122898 90772
rect 167730 90760 167736 90772
rect 122892 90732 167736 90760
rect 122892 90720 122898 90732
rect 167730 90720 167736 90732
rect 167788 90720 167794 90772
rect 151722 90652 151728 90704
rect 151780 90692 151786 90704
rect 184198 90692 184204 90704
rect 151780 90664 184204 90692
rect 151780 90652 151786 90664
rect 184198 90652 184204 90664
rect 184256 90652 184262 90704
rect 309686 90380 309692 90432
rect 309744 90420 309750 90432
rect 320174 90420 320180 90432
rect 309744 90392 320180 90420
rect 309744 90380 309750 90392
rect 320174 90380 320180 90392
rect 320232 90380 320238 90432
rect 308582 90312 308588 90364
rect 308640 90352 308646 90364
rect 328454 90352 328460 90364
rect 308640 90324 328460 90352
rect 308640 90312 308646 90324
rect 328454 90312 328460 90324
rect 328512 90312 328518 90364
rect 89070 89632 89076 89684
rect 89128 89672 89134 89684
rect 209130 89672 209136 89684
rect 89128 89644 209136 89672
rect 89128 89632 89134 89644
rect 209130 89632 209136 89644
rect 209188 89632 209194 89684
rect 123938 89564 123944 89616
rect 123996 89604 124002 89616
rect 213178 89604 213184 89616
rect 123996 89576 213184 89604
rect 123996 89564 124002 89576
rect 213178 89564 213184 89576
rect 213236 89564 213242 89616
rect 112346 89496 112352 89548
rect 112404 89536 112410 89548
rect 182910 89536 182916 89548
rect 112404 89508 182916 89536
rect 112404 89496 112410 89508
rect 182910 89496 182916 89508
rect 182968 89496 182974 89548
rect 104526 89428 104532 89480
rect 104584 89468 104590 89480
rect 170582 89468 170588 89480
rect 104584 89440 170588 89468
rect 104584 89428 104590 89440
rect 170582 89428 170588 89440
rect 170640 89428 170646 89480
rect 106918 89360 106924 89412
rect 106976 89400 106982 89412
rect 173158 89400 173164 89412
rect 106976 89372 173164 89400
rect 106976 89360 106982 89372
rect 173158 89360 173164 89372
rect 173216 89360 173222 89412
rect 126606 89292 126612 89344
rect 126664 89332 126670 89344
rect 166350 89332 166356 89344
rect 126664 89304 166356 89332
rect 126664 89292 126670 89304
rect 166350 89292 166356 89304
rect 166408 89292 166414 89344
rect 91002 88272 91008 88324
rect 91060 88312 91066 88324
rect 212074 88312 212080 88324
rect 91060 88284 212080 88312
rect 91060 88272 91066 88284
rect 212074 88272 212080 88284
rect 212132 88272 212138 88324
rect 106642 88204 106648 88256
rect 106700 88244 106706 88256
rect 203610 88244 203616 88256
rect 106700 88216 203616 88244
rect 106700 88204 106706 88216
rect 203610 88204 203616 88216
rect 203668 88204 203674 88256
rect 87414 88136 87420 88188
rect 87472 88176 87478 88188
rect 164878 88176 164884 88188
rect 87472 88148 164884 88176
rect 87472 88136 87478 88148
rect 164878 88136 164884 88148
rect 164936 88136 164942 88188
rect 110138 88068 110144 88120
rect 110196 88108 110202 88120
rect 167822 88108 167828 88120
rect 110196 88080 167828 88108
rect 110196 88068 110202 88080
rect 167822 88068 167828 88080
rect 167880 88068 167886 88120
rect 135898 88000 135904 88052
rect 135956 88040 135962 88052
rect 185670 88040 185676 88052
rect 135956 88012 185676 88040
rect 135956 88000 135962 88012
rect 185670 88000 185676 88012
rect 185728 88000 185734 88052
rect 121086 87932 121092 87984
rect 121144 87972 121150 87984
rect 170490 87972 170496 87984
rect 121144 87944 170496 87972
rect 121144 87932 121150 87944
rect 170490 87932 170496 87944
rect 170548 87932 170554 87984
rect 300118 87660 300124 87712
rect 300176 87700 300182 87712
rect 324314 87700 324320 87712
rect 300176 87672 324320 87700
rect 300176 87660 300182 87672
rect 324314 87660 324320 87672
rect 324372 87660 324378 87712
rect 3510 87592 3516 87644
rect 3568 87632 3574 87644
rect 21358 87632 21364 87644
rect 3568 87604 21364 87632
rect 3568 87592 3574 87604
rect 21358 87592 21364 87604
rect 21416 87592 21422 87644
rect 185578 87592 185584 87644
rect 185636 87632 185642 87644
rect 307294 87632 307300 87644
rect 185636 87604 307300 87632
rect 185636 87592 185642 87604
rect 307294 87592 307300 87604
rect 307352 87592 307358 87644
rect 63402 86912 63408 86964
rect 63460 86952 63466 86964
rect 206370 86952 206376 86964
rect 63460 86924 206376 86952
rect 63460 86912 63466 86924
rect 206370 86912 206376 86924
rect 206428 86912 206434 86964
rect 274082 86912 274088 86964
rect 274140 86952 274146 86964
rect 580166 86952 580172 86964
rect 274140 86924 580172 86952
rect 274140 86912 274146 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 99926 86844 99932 86896
rect 99984 86884 99990 86896
rect 200758 86884 200764 86896
rect 99984 86856 200764 86884
rect 99984 86844 99990 86856
rect 200758 86844 200764 86856
rect 200816 86844 200822 86896
rect 117130 86776 117136 86828
rect 117188 86816 117194 86828
rect 213270 86816 213276 86828
rect 117188 86788 213276 86816
rect 117188 86776 117194 86788
rect 213270 86776 213276 86788
rect 213328 86776 213334 86828
rect 102962 86708 102968 86760
rect 103020 86748 103026 86760
rect 177390 86748 177396 86760
rect 103020 86720 177396 86748
rect 103020 86708 103026 86720
rect 177390 86708 177396 86720
rect 177448 86708 177454 86760
rect 122374 86640 122380 86692
rect 122432 86680 122438 86692
rect 193858 86680 193864 86692
rect 122432 86652 193864 86680
rect 122432 86640 122438 86652
rect 193858 86640 193864 86652
rect 193916 86640 193922 86692
rect 252554 86232 252560 86284
rect 252612 86272 252618 86284
rect 291930 86272 291936 86284
rect 252612 86244 291936 86272
rect 252612 86232 252618 86244
rect 291930 86232 291936 86244
rect 291988 86232 291994 86284
rect 67634 85484 67640 85536
rect 67692 85524 67698 85536
rect 214834 85524 214840 85536
rect 67692 85496 214840 85524
rect 67692 85484 67698 85496
rect 214834 85484 214840 85496
rect 214892 85484 214898 85536
rect 85022 85416 85028 85468
rect 85080 85456 85086 85468
rect 173434 85456 173440 85468
rect 85080 85428 173440 85456
rect 85080 85416 85086 85428
rect 173434 85416 173440 85428
rect 173492 85416 173498 85468
rect 96522 85348 96528 85400
rect 96580 85388 96586 85400
rect 167914 85388 167920 85400
rect 96580 85360 167920 85388
rect 96580 85348 96586 85360
rect 167914 85348 167920 85360
rect 167972 85348 167978 85400
rect 118234 85280 118240 85332
rect 118292 85320 118298 85332
rect 188430 85320 188436 85332
rect 118292 85292 188436 85320
rect 118292 85280 118298 85292
rect 188430 85280 188436 85292
rect 188488 85280 188494 85332
rect 135070 85212 135076 85264
rect 135128 85252 135134 85264
rect 203518 85252 203524 85264
rect 135128 85224 203524 85252
rect 135128 85212 135134 85224
rect 203518 85212 203524 85224
rect 203576 85212 203582 85264
rect 116762 85144 116768 85196
rect 116820 85184 116826 85196
rect 169110 85184 169116 85196
rect 116820 85156 169116 85184
rect 116820 85144 116826 85156
rect 169110 85144 169116 85156
rect 169168 85144 169174 85196
rect 238754 84872 238760 84924
rect 238812 84912 238818 84924
rect 295426 84912 295432 84924
rect 238812 84884 295432 84912
rect 238812 84872 238818 84884
rect 295426 84872 295432 84884
rect 295484 84872 295490 84924
rect 179230 84804 179236 84856
rect 179288 84844 179294 84856
rect 267826 84844 267832 84856
rect 179288 84816 267832 84844
rect 179288 84804 179294 84816
rect 267826 84804 267832 84816
rect 267884 84804 267890 84856
rect 64690 84124 64696 84176
rect 64748 84164 64754 84176
rect 193950 84164 193956 84176
rect 64748 84136 193956 84164
rect 64748 84124 64754 84136
rect 193950 84124 193956 84136
rect 194008 84124 194014 84176
rect 112438 84056 112444 84108
rect 112496 84096 112502 84108
rect 214650 84096 214656 84108
rect 112496 84068 214656 84096
rect 112496 84056 112502 84068
rect 214650 84056 214656 84068
rect 214708 84056 214714 84108
rect 119982 83988 119988 84040
rect 120040 84028 120046 84040
rect 210510 84028 210516 84040
rect 120040 84000 210516 84028
rect 120040 83988 120046 84000
rect 210510 83988 210516 84000
rect 210568 83988 210574 84040
rect 106182 83920 106188 83972
rect 106240 83960 106246 83972
rect 173250 83960 173256 83972
rect 106240 83932 173256 83960
rect 106240 83920 106246 83932
rect 173250 83920 173256 83932
rect 173308 83920 173314 83972
rect 129642 83852 129648 83904
rect 129700 83892 129706 83904
rect 167638 83892 167644 83904
rect 129700 83864 167644 83892
rect 129700 83852 129706 83864
rect 167638 83852 167644 83864
rect 167696 83852 167702 83904
rect 285766 83512 285772 83564
rect 285824 83552 285830 83564
rect 293034 83552 293040 83564
rect 285824 83524 293040 83552
rect 285824 83512 285830 83524
rect 293034 83512 293040 83524
rect 293092 83512 293098 83564
rect 176470 83444 176476 83496
rect 176528 83484 176534 83496
rect 313274 83484 313280 83496
rect 176528 83456 313280 83484
rect 176528 83444 176534 83456
rect 313274 83444 313280 83456
rect 313332 83444 313338 83496
rect 100662 82764 100668 82816
rect 100720 82804 100726 82816
rect 189902 82804 189908 82816
rect 100720 82776 189908 82804
rect 100720 82764 100726 82776
rect 189902 82764 189908 82776
rect 189960 82764 189966 82816
rect 126882 82696 126888 82748
rect 126940 82736 126946 82748
rect 209038 82736 209044 82748
rect 126940 82708 209044 82736
rect 126940 82696 126946 82708
rect 209038 82696 209044 82708
rect 209096 82696 209102 82748
rect 115750 82628 115756 82680
rect 115808 82668 115814 82680
rect 196802 82668 196808 82680
rect 115808 82640 196808 82668
rect 115808 82628 115814 82640
rect 196802 82628 196808 82640
rect 196860 82628 196866 82680
rect 86770 82560 86776 82612
rect 86828 82600 86834 82612
rect 166534 82600 166540 82612
rect 86828 82572 166540 82600
rect 86828 82560 86834 82572
rect 166534 82560 166540 82572
rect 166592 82560 166598 82612
rect 103422 82492 103428 82544
rect 103480 82532 103486 82544
rect 171870 82532 171876 82544
rect 103480 82504 171876 82532
rect 103480 82492 103486 82504
rect 171870 82492 171876 82504
rect 171928 82492 171934 82544
rect 198090 82220 198096 82272
rect 198148 82260 198154 82272
rect 260098 82260 260104 82272
rect 198148 82232 260104 82260
rect 198148 82220 198154 82232
rect 260098 82220 260104 82232
rect 260156 82220 260162 82272
rect 216030 82152 216036 82204
rect 216088 82192 216094 82204
rect 327074 82192 327080 82204
rect 216088 82164 327080 82192
rect 216088 82152 216094 82164
rect 327074 82152 327080 82164
rect 327132 82152 327138 82204
rect 191098 82084 191104 82136
rect 191156 82124 191162 82136
rect 323578 82124 323584 82136
rect 191156 82096 323584 82124
rect 191156 82084 191162 82096
rect 323578 82084 323584 82096
rect 323636 82084 323642 82136
rect 45186 81336 45192 81388
rect 45244 81376 45250 81388
rect 322934 81376 322940 81388
rect 45244 81348 322940 81376
rect 45244 81336 45250 81348
rect 322934 81336 322940 81348
rect 322992 81336 322998 81388
rect 92382 81268 92388 81320
rect 92440 81308 92446 81320
rect 192754 81308 192760 81320
rect 92440 81280 192760 81308
rect 92440 81268 92446 81280
rect 192754 81268 192760 81280
rect 192812 81268 192818 81320
rect 95050 81200 95056 81252
rect 95108 81240 95114 81252
rect 188522 81240 188528 81252
rect 95108 81212 188528 81240
rect 95108 81200 95114 81212
rect 188522 81200 188528 81212
rect 188580 81200 188586 81252
rect 131022 81132 131028 81184
rect 131080 81172 131086 81184
rect 211890 81172 211896 81184
rect 131080 81144 211896 81172
rect 131080 81132 131086 81144
rect 211890 81132 211896 81144
rect 211948 81132 211954 81184
rect 120810 81064 120816 81116
rect 120868 81104 120874 81116
rect 187142 81104 187148 81116
rect 120868 81076 187148 81104
rect 120868 81064 120874 81076
rect 187142 81064 187148 81076
rect 187200 81064 187206 81116
rect 35802 79976 35808 80028
rect 35860 80016 35866 80028
rect 321830 80016 321836 80028
rect 35860 79988 321836 80016
rect 35860 79976 35866 79988
rect 321830 79976 321836 79988
rect 321888 79976 321894 80028
rect 102042 79908 102048 79960
rect 102100 79948 102106 79960
rect 188338 79948 188344 79960
rect 102100 79920 188344 79948
rect 102100 79908 102106 79920
rect 188338 79908 188344 79920
rect 188396 79908 188402 79960
rect 120718 79840 120724 79892
rect 120776 79880 120782 79892
rect 205082 79880 205088 79892
rect 120776 79852 205088 79880
rect 120776 79840 120782 79852
rect 205082 79840 205088 79852
rect 205140 79840 205146 79892
rect 97810 79772 97816 79824
rect 97868 79812 97874 79824
rect 178678 79812 178684 79824
rect 97868 79784 178684 79812
rect 97868 79772 97874 79784
rect 178678 79772 178684 79784
rect 178736 79772 178742 79824
rect 99098 79704 99104 79756
rect 99156 79744 99162 79756
rect 171962 79744 171968 79756
rect 99156 79716 171968 79744
rect 99156 79704 99162 79716
rect 171962 79704 171968 79716
rect 172020 79704 172026 79756
rect 39850 78616 39856 78668
rect 39908 78656 39914 78668
rect 318058 78656 318064 78668
rect 39908 78628 318064 78656
rect 39908 78616 39914 78628
rect 318058 78616 318064 78628
rect 318116 78616 318122 78668
rect 97902 78548 97908 78600
rect 97960 78588 97966 78600
rect 189810 78588 189816 78600
rect 97960 78560 189816 78588
rect 97960 78548 97966 78560
rect 189810 78548 189816 78560
rect 189868 78548 189874 78600
rect 125502 78480 125508 78532
rect 125560 78520 125566 78532
rect 211982 78520 211988 78532
rect 125560 78492 211988 78520
rect 125560 78480 125566 78492
rect 211982 78480 211988 78492
rect 212040 78480 212046 78532
rect 118602 78412 118608 78464
rect 118660 78452 118666 78464
rect 192662 78452 192668 78464
rect 118660 78424 192668 78452
rect 118660 78412 118666 78424
rect 192662 78412 192668 78424
rect 192720 78412 192726 78464
rect 99282 77188 99288 77240
rect 99340 77228 99346 77240
rect 184290 77228 184296 77240
rect 99340 77200 184296 77228
rect 99340 77188 99346 77200
rect 184290 77188 184296 77200
rect 184348 77188 184354 77240
rect 114462 77120 114468 77172
rect 114520 77160 114526 77172
rect 169018 77160 169024 77172
rect 114520 77132 169024 77160
rect 114520 77120 114526 77132
rect 169018 77120 169024 77132
rect 169076 77120 169082 77172
rect 115934 76576 115940 76628
rect 115992 76616 115998 76628
rect 301774 76616 301780 76628
rect 115992 76588 301780 76616
rect 115992 76576 115998 76588
rect 301774 76576 301780 76588
rect 301832 76576 301838 76628
rect 80054 76508 80060 76560
rect 80112 76548 80118 76560
rect 304534 76548 304540 76560
rect 80112 76520 304540 76548
rect 80112 76508 80118 76520
rect 304534 76508 304540 76520
rect 304592 76508 304598 76560
rect 308398 76508 308404 76560
rect 308456 76548 308462 76560
rect 316126 76548 316132 76560
rect 308456 76520 316132 76548
rect 308456 76508 308462 76520
rect 316126 76508 316132 76520
rect 316184 76508 316190 76560
rect 93762 75828 93768 75880
rect 93820 75868 93826 75880
rect 174630 75868 174636 75880
rect 93820 75840 174636 75868
rect 93820 75828 93826 75840
rect 174630 75828 174636 75840
rect 174688 75828 174694 75880
rect 111702 75760 111708 75812
rect 111760 75800 111766 75812
rect 185762 75800 185768 75812
rect 111760 75772 185768 75800
rect 111760 75760 111766 75772
rect 185762 75760 185768 75772
rect 185820 75760 185826 75812
rect 184934 75216 184940 75268
rect 184992 75256 184998 75268
rect 315298 75256 315304 75268
rect 184992 75228 315304 75256
rect 184992 75216 184998 75228
rect 315298 75216 315304 75228
rect 315356 75216 315362 75268
rect 97994 75148 98000 75200
rect 98052 75188 98058 75200
rect 285122 75188 285128 75200
rect 98052 75160 285128 75188
rect 98052 75148 98058 75160
rect 285122 75148 285128 75160
rect 285180 75148 285186 75200
rect 127618 74468 127624 74520
rect 127676 74508 127682 74520
rect 207750 74508 207756 74520
rect 127676 74480 207756 74508
rect 127676 74468 127682 74480
rect 207750 74468 207756 74480
rect 207808 74468 207814 74520
rect 81434 73856 81440 73908
rect 81492 73896 81498 73908
rect 305730 73896 305736 73908
rect 81492 73868 305736 73896
rect 81492 73856 81498 73868
rect 305730 73856 305736 73868
rect 305788 73856 305794 73908
rect 6914 73788 6920 73840
rect 6972 73828 6978 73840
rect 293402 73828 293408 73840
rect 6972 73800 293408 73828
rect 6972 73788 6978 73800
rect 293402 73788 293408 73800
rect 293460 73788 293466 73840
rect 309870 73652 309876 73704
rect 309928 73692 309934 73704
rect 317414 73692 317420 73704
rect 309928 73664 317420 73692
rect 309928 73652 309934 73664
rect 317414 73652 317420 73664
rect 317472 73652 317478 73704
rect 356698 73108 356704 73160
rect 356756 73148 356762 73160
rect 580166 73148 580172 73160
rect 356756 73120 580172 73148
rect 356756 73108 356762 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 85574 72496 85580 72548
rect 85632 72536 85638 72548
rect 279510 72536 279516 72548
rect 85632 72508 279516 72536
rect 85632 72496 85638 72508
rect 279510 72496 279516 72508
rect 279568 72496 279574 72548
rect 46934 72428 46940 72480
rect 46992 72468 46998 72480
rect 296162 72468 296168 72480
rect 46992 72440 296168 72468
rect 46992 72428 46998 72440
rect 296162 72428 296168 72440
rect 296220 72428 296226 72480
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 43438 71720 43444 71732
rect 3476 71692 43444 71720
rect 3476 71680 3482 71692
rect 43438 71680 43444 71692
rect 43496 71680 43502 71732
rect 113174 71136 113180 71188
rect 113232 71176 113238 71188
rect 297542 71176 297548 71188
rect 113232 71148 297548 71176
rect 113232 71136 113238 71148
rect 297542 71136 297548 71148
rect 297600 71136 297606 71188
rect 44174 71068 44180 71120
rect 44232 71108 44238 71120
rect 261662 71108 261668 71120
rect 44232 71080 261668 71108
rect 44232 71068 44238 71080
rect 261662 71068 261668 71080
rect 261720 71068 261726 71120
rect 37274 71000 37280 71052
rect 37332 71040 37338 71052
rect 304442 71040 304448 71052
rect 37332 71012 304448 71040
rect 37332 71000 37338 71012
rect 304442 71000 304448 71012
rect 304500 71000 304506 71052
rect 51074 69640 51080 69692
rect 51132 69680 51138 69692
rect 294874 69680 294880 69692
rect 51132 69652 294880 69680
rect 51132 69640 51138 69652
rect 294874 69640 294880 69652
rect 294932 69640 294938 69692
rect 92474 68348 92480 68400
rect 92532 68388 92538 68400
rect 294690 68388 294696 68400
rect 92532 68360 294696 68388
rect 92532 68348 92538 68360
rect 294690 68348 294696 68360
rect 294748 68348 294754 68400
rect 57974 68280 57980 68332
rect 58032 68320 58038 68332
rect 303154 68320 303160 68332
rect 58032 68292 303160 68320
rect 58032 68280 58038 68292
rect 303154 68280 303160 68292
rect 303212 68280 303218 68332
rect 99374 66920 99380 66972
rect 99432 66960 99438 66972
rect 278314 66960 278320 66972
rect 99432 66932 278320 66960
rect 99432 66920 99438 66932
rect 278314 66920 278320 66932
rect 278372 66920 278378 66972
rect 64874 66852 64880 66904
rect 64932 66892 64938 66904
rect 296070 66892 296076 66904
rect 64932 66864 296076 66892
rect 64932 66852 64938 66864
rect 296070 66852 296076 66864
rect 296128 66852 296134 66904
rect 106274 65560 106280 65612
rect 106332 65600 106338 65612
rect 266998 65600 267004 65612
rect 106332 65572 267004 65600
rect 106332 65560 106338 65572
rect 266998 65560 267004 65572
rect 267056 65560 267062 65612
rect 69014 65492 69020 65544
rect 69072 65532 69078 65544
rect 305914 65532 305920 65544
rect 69072 65504 305920 65532
rect 69072 65492 69078 65504
rect 305914 65492 305920 65504
rect 305972 65492 305978 65544
rect 71774 64200 71780 64252
rect 71832 64240 71838 64252
rect 261570 64240 261576 64252
rect 71832 64212 261576 64240
rect 71832 64200 71838 64212
rect 261570 64200 261576 64212
rect 261628 64200 261634 64252
rect 34514 64132 34520 64184
rect 34572 64172 34578 64184
rect 297634 64172 297640 64184
rect 34572 64144 297640 64172
rect 34572 64132 34578 64144
rect 297634 64132 297640 64144
rect 297692 64132 297698 64184
rect 110414 62840 110420 62892
rect 110472 62880 110478 62892
rect 250622 62880 250628 62892
rect 110472 62852 250628 62880
rect 110472 62840 110478 62852
rect 250622 62840 250628 62852
rect 250680 62840 250686 62892
rect 117314 62772 117320 62824
rect 117372 62812 117378 62824
rect 290550 62812 290556 62824
rect 117372 62784 290556 62812
rect 117372 62772 117378 62784
rect 290550 62772 290556 62784
rect 290608 62772 290614 62824
rect 82814 61412 82820 61464
rect 82872 61452 82878 61464
rect 267090 61452 267096 61464
rect 82872 61424 267096 61452
rect 82872 61412 82878 61424
rect 267090 61412 267096 61424
rect 267148 61412 267154 61464
rect 67634 61344 67640 61396
rect 67692 61384 67698 61396
rect 301590 61384 301596 61396
rect 67692 61356 301596 61384
rect 67692 61344 67698 61356
rect 301590 61344 301596 61356
rect 301648 61344 301654 61396
rect 359458 60664 359464 60716
rect 359516 60704 359522 60716
rect 580166 60704 580172 60716
rect 359516 60676 580172 60704
rect 359516 60664 359522 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 85666 59984 85672 60036
rect 85724 60024 85730 60036
rect 303062 60024 303068 60036
rect 85724 59996 303068 60024
rect 85724 59984 85730 59996
rect 303062 59984 303068 59996
rect 303120 59984 303126 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 58618 59344 58624 59356
rect 3108 59316 58624 59344
rect 3108 59304 3114 59316
rect 58618 59304 58624 59316
rect 58676 59304 58682 59356
rect 120074 58692 120080 58744
rect 120132 58732 120138 58744
rect 272518 58732 272524 58744
rect 120132 58704 272524 58732
rect 120132 58692 120138 58704
rect 272518 58692 272524 58704
rect 272576 58692 272582 58744
rect 89714 58624 89720 58676
rect 89772 58664 89778 58676
rect 300394 58664 300400 58676
rect 89772 58636 300400 58664
rect 89772 58624 89778 58636
rect 300394 58624 300400 58636
rect 300452 58624 300458 58676
rect 74534 57264 74540 57316
rect 74592 57304 74598 57316
rect 282270 57304 282276 57316
rect 74592 57276 282276 57304
rect 74592 57264 74598 57276
rect 282270 57264 282276 57276
rect 282328 57264 282334 57316
rect 93854 57196 93860 57248
rect 93912 57236 93918 57248
rect 305822 57236 305828 57248
rect 93912 57208 305828 57236
rect 93912 57196 93918 57208
rect 305822 57196 305828 57208
rect 305880 57196 305886 57248
rect 96614 55904 96620 55956
rect 96672 55944 96678 55956
rect 271230 55944 271236 55956
rect 96672 55916 271236 55944
rect 96672 55904 96678 55916
rect 271230 55904 271236 55916
rect 271288 55904 271294 55956
rect 70394 55836 70400 55888
rect 70452 55876 70458 55888
rect 280982 55876 280988 55888
rect 70452 55848 280988 55876
rect 70452 55836 70458 55848
rect 280982 55836 280988 55848
rect 281040 55836 281046 55888
rect 100754 54544 100760 54596
rect 100812 54584 100818 54596
rect 299014 54584 299020 54596
rect 100812 54556 299020 54584
rect 100812 54544 100818 54556
rect 299014 54544 299020 54556
rect 299072 54544 299078 54596
rect 63494 54476 63500 54528
rect 63552 54516 63558 54528
rect 283834 54516 283840 54528
rect 63552 54488 283840 54516
rect 63552 54476 63558 54488
rect 283834 54476 283840 54488
rect 283892 54476 283898 54528
rect 103514 53116 103520 53168
rect 103572 53156 103578 53168
rect 304350 53156 304356 53168
rect 103572 53128 304356 53156
rect 103572 53116 103578 53128
rect 304350 53116 304356 53128
rect 304408 53116 304414 53168
rect 60734 53048 60740 53100
rect 60792 53088 60798 53100
rect 285030 53088 285036 53100
rect 60792 53060 285036 53088
rect 60792 53048 60798 53060
rect 285030 53048 285036 53060
rect 285088 53048 285094 53100
rect 107654 51756 107660 51808
rect 107712 51796 107718 51808
rect 275370 51796 275376 51808
rect 107712 51768 275376 51796
rect 107712 51756 107718 51768
rect 275370 51756 275376 51768
rect 275428 51756 275434 51808
rect 4154 51688 4160 51740
rect 4212 51728 4218 51740
rect 307202 51728 307208 51740
rect 4212 51700 307208 51728
rect 4212 51688 4218 51700
rect 307202 51688 307208 51700
rect 307260 51688 307266 51740
rect 84194 50396 84200 50448
rect 84252 50436 84258 50448
rect 298922 50436 298928 50448
rect 84252 50408 298928 50436
rect 84252 50396 84258 50408
rect 298922 50396 298928 50408
rect 298980 50396 298986 50448
rect 44266 50328 44272 50380
rect 44324 50368 44330 50380
rect 262950 50368 262956 50380
rect 44324 50340 262956 50368
rect 44324 50328 44330 50340
rect 262950 50328 262956 50340
rect 263008 50328 263014 50380
rect 102134 49036 102140 49088
rect 102192 49076 102198 49088
rect 250438 49076 250444 49088
rect 102192 49048 250444 49076
rect 102192 49036 102198 49048
rect 250438 49036 250444 49048
rect 250496 49036 250502 49088
rect 124214 48968 124220 49020
rect 124272 49008 124278 49020
rect 280890 49008 280896 49020
rect 124272 48980 280896 49008
rect 124272 48968 124278 48980
rect 280890 48968 280896 48980
rect 280948 48968 280954 49020
rect 30374 47608 30380 47660
rect 30432 47648 30438 47660
rect 268470 47648 268476 47660
rect 30432 47620 268476 47648
rect 30432 47608 30438 47620
rect 268470 47608 268476 47620
rect 268528 47608 268534 47660
rect 49694 47540 49700 47592
rect 49752 47580 49758 47592
rect 307110 47580 307116 47592
rect 49752 47552 307116 47580
rect 49752 47540 49758 47552
rect 307110 47540 307116 47552
rect 307168 47540 307174 47592
rect 353938 46860 353944 46912
rect 353996 46900 354002 46912
rect 580166 46900 580172 46912
rect 353996 46872 580172 46900
rect 353996 46860 354002 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 35986 46248 35992 46300
rect 36044 46288 36050 46300
rect 287790 46288 287796 46300
rect 36044 46260 287796 46288
rect 36044 46248 36050 46260
rect 287790 46248 287796 46260
rect 287848 46248 287854 46300
rect 20714 46180 20720 46232
rect 20772 46220 20778 46232
rect 289262 46220 289268 46232
rect 20772 46192 289268 46220
rect 20772 46180 20778 46192
rect 289262 46180 289268 46192
rect 289320 46180 289326 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 18598 45540 18604 45552
rect 3476 45512 18604 45540
rect 3476 45500 3482 45512
rect 18598 45500 18604 45512
rect 18656 45500 18662 45552
rect 19334 44888 19340 44940
rect 19392 44928 19398 44940
rect 260190 44928 260196 44940
rect 19392 44900 260196 44928
rect 19392 44888 19398 44900
rect 260190 44888 260196 44900
rect 260248 44888 260254 44940
rect 40034 44820 40040 44872
rect 40092 44860 40098 44872
rect 294782 44860 294788 44872
rect 40092 44832 294788 44860
rect 40092 44820 40098 44832
rect 294782 44820 294788 44832
rect 294840 44820 294846 44872
rect 102226 43460 102232 43512
rect 102284 43500 102290 43512
rect 287882 43500 287888 43512
rect 102284 43472 287888 43500
rect 102284 43460 102290 43472
rect 287882 43460 287888 43472
rect 287940 43460 287946 43512
rect 38654 43392 38660 43444
rect 38712 43432 38718 43444
rect 269850 43432 269856 43444
rect 38712 43404 269856 43432
rect 38712 43392 38718 43404
rect 269850 43392 269856 43404
rect 269908 43392 269914 43444
rect 118694 42100 118700 42152
rect 118752 42140 118758 42152
rect 300302 42140 300308 42152
rect 118752 42112 300308 42140
rect 118752 42100 118758 42112
rect 300302 42100 300308 42112
rect 300360 42100 300366 42152
rect 41414 42032 41420 42084
rect 41472 42072 41478 42084
rect 282362 42072 282368 42084
rect 41472 42044 282368 42072
rect 41472 42032 41478 42044
rect 282362 42032 282368 42044
rect 282420 42032 282426 42084
rect 110506 40740 110512 40792
rect 110564 40780 110570 40792
rect 304258 40780 304264 40792
rect 110564 40752 304264 40780
rect 110564 40740 110570 40752
rect 304258 40740 304264 40752
rect 304316 40740 304322 40792
rect 9674 40672 9680 40724
rect 9732 40712 9738 40724
rect 289170 40712 289176 40724
rect 9732 40684 289176 40712
rect 9732 40672 9738 40684
rect 289170 40672 289176 40684
rect 289228 40672 289234 40724
rect 42794 39380 42800 39432
rect 42852 39420 42858 39432
rect 278222 39420 278228 39432
rect 42852 39392 278228 39420
rect 42852 39380 42858 39392
rect 278222 39380 278228 39392
rect 278280 39380 278286 39432
rect 11054 39312 11060 39364
rect 11112 39352 11118 39364
rect 274174 39352 274180 39364
rect 11112 39324 274180 39352
rect 11112 39312 11118 39324
rect 274174 39312 274180 39324
rect 274232 39312 274238 39364
rect 45554 37884 45560 37936
rect 45612 37924 45618 37936
rect 273990 37924 273996 37936
rect 45612 37896 273996 37924
rect 45612 37884 45618 37896
rect 273990 37884 273996 37896
rect 274048 37884 274054 37936
rect 78674 36592 78680 36644
rect 78732 36632 78738 36644
rect 301682 36632 301688 36644
rect 78732 36604 301688 36632
rect 78732 36592 78738 36604
rect 301682 36592 301688 36604
rect 301740 36592 301746 36644
rect 19426 36524 19432 36576
rect 19484 36564 19490 36576
rect 271138 36564 271144 36576
rect 19484 36536 271144 36564
rect 19484 36524 19490 36536
rect 271138 36524 271144 36536
rect 271196 36524 271202 36576
rect 128354 35232 128360 35284
rect 128412 35272 128418 35284
rect 216674 35272 216680 35284
rect 128412 35244 216680 35272
rect 128412 35232 128418 35244
rect 216674 35232 216680 35244
rect 216732 35232 216738 35284
rect 238018 35232 238024 35284
rect 238076 35272 238082 35284
rect 251358 35272 251364 35284
rect 238076 35244 251364 35272
rect 238076 35232 238082 35244
rect 251358 35232 251364 35244
rect 251416 35232 251422 35284
rect 12434 35164 12440 35216
rect 12492 35204 12498 35216
rect 294598 35204 294604 35216
rect 12492 35176 294604 35204
rect 12492 35164 12498 35176
rect 294598 35164 294604 35176
rect 294656 35164 294662 35216
rect 53834 33804 53840 33856
rect 53892 33844 53898 33856
rect 293310 33844 293316 33856
rect 53892 33816 293316 33844
rect 53892 33804 53898 33816
rect 293310 33804 293316 33816
rect 293368 33804 293374 33856
rect 31754 33736 31760 33788
rect 31812 33776 31818 33788
rect 286318 33776 286324 33788
rect 31812 33748 286324 33776
rect 31812 33736 31818 33748
rect 286318 33736 286324 33748
rect 286376 33736 286382 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 46198 33096 46204 33108
rect 3568 33068 46204 33096
rect 3568 33056 3574 33068
rect 46198 33056 46204 33068
rect 46256 33056 46262 33108
rect 345658 33056 345664 33108
rect 345716 33096 345722 33108
rect 579890 33096 579896 33108
rect 345716 33068 579896 33096
rect 345716 33056 345722 33068
rect 579890 33056 579896 33068
rect 579948 33056 579954 33108
rect 180794 32512 180800 32564
rect 180852 32552 180858 32564
rect 261570 32552 261576 32564
rect 180852 32524 261576 32552
rect 180852 32512 180858 32524
rect 261570 32512 261576 32524
rect 261628 32512 261634 32564
rect 201494 32444 201500 32496
rect 201552 32484 201558 32496
rect 343634 32484 343640 32496
rect 201552 32456 343640 32484
rect 201552 32444 201558 32456
rect 343634 32444 343640 32456
rect 343692 32444 343698 32496
rect 93946 32376 93952 32428
rect 94004 32416 94010 32428
rect 300210 32416 300216 32428
rect 94004 32388 300216 32416
rect 94004 32376 94010 32388
rect 300210 32376 300216 32388
rect 300268 32376 300274 32428
rect 200114 31152 200120 31204
rect 200172 31192 200178 31204
rect 311894 31192 311900 31204
rect 200172 31164 311900 31192
rect 200172 31152 200178 31164
rect 311894 31152 311900 31164
rect 311952 31152 311958 31204
rect 104894 31084 104900 31136
rect 104952 31124 104958 31136
rect 290458 31124 290464 31136
rect 104952 31096 290464 31124
rect 104952 31084 104958 31096
rect 290458 31084 290464 31096
rect 290516 31084 290522 31136
rect 75914 31016 75920 31068
rect 75972 31056 75978 31068
rect 276658 31056 276664 31068
rect 75972 31028 276664 31056
rect 75972 31016 75978 31028
rect 276658 31016 276664 31028
rect 276716 31016 276722 31068
rect 73154 29656 73160 29708
rect 73212 29696 73218 29708
rect 269758 29696 269764 29708
rect 73212 29668 269764 29696
rect 73212 29656 73218 29668
rect 269758 29656 269764 29668
rect 269816 29656 269822 29708
rect 17954 29588 17960 29640
rect 18012 29628 18018 29640
rect 284938 29628 284944 29640
rect 18012 29600 284944 29628
rect 18012 29588 18018 29600
rect 284938 29588 284944 29600
rect 284996 29588 285002 29640
rect 86954 28296 86960 28348
rect 87012 28336 87018 28348
rect 261478 28336 261484 28348
rect 87012 28308 261484 28336
rect 87012 28296 87018 28308
rect 261478 28296 261484 28308
rect 261536 28296 261542 28348
rect 22094 28228 22100 28280
rect 22152 28268 22158 28280
rect 307018 28268 307024 28280
rect 22152 28240 307024 28268
rect 22152 28228 22158 28240
rect 307018 28228 307024 28240
rect 307076 28228 307082 28280
rect 297358 27548 297364 27600
rect 297416 27588 297422 27600
rect 299474 27588 299480 27600
rect 297416 27560 299480 27588
rect 297416 27548 297422 27560
rect 299474 27548 299480 27560
rect 299532 27548 299538 27600
rect 179322 26936 179328 26988
rect 179380 26976 179386 26988
rect 273254 26976 273260 26988
rect 179380 26948 273260 26976
rect 179380 26936 179386 26948
rect 273254 26936 273260 26948
rect 273312 26936 273318 26988
rect 26234 26868 26240 26920
rect 26292 26908 26298 26920
rect 250530 26908 250536 26920
rect 26292 26880 250536 26908
rect 26292 26868 26298 26880
rect 250530 26868 250536 26880
rect 250588 26868 250594 26920
rect 210418 25644 210424 25696
rect 210476 25684 210482 25696
rect 324406 25684 324412 25696
rect 210476 25656 324412 25684
rect 210476 25644 210482 25656
rect 324406 25644 324412 25656
rect 324464 25644 324470 25696
rect 176562 25576 176568 25628
rect 176620 25616 176626 25628
rect 296714 25616 296720 25628
rect 176620 25588 296720 25616
rect 176620 25576 176626 25588
rect 296714 25576 296720 25588
rect 296772 25576 296778 25628
rect 77294 25508 77300 25560
rect 77352 25548 77358 25560
rect 273898 25548 273904 25560
rect 77352 25520 273904 25548
rect 77352 25508 77358 25520
rect 273898 25508 273904 25520
rect 273956 25508 273962 25560
rect 62114 24148 62120 24200
rect 62172 24188 62178 24200
rect 302970 24188 302976 24200
rect 62172 24160 302976 24188
rect 62172 24148 62178 24160
rect 302970 24148 302976 24160
rect 303028 24148 303034 24200
rect 2866 24080 2872 24132
rect 2924 24120 2930 24132
rect 262858 24120 262864 24132
rect 2924 24092 262864 24120
rect 2924 24080 2930 24092
rect 262858 24080 262864 24092
rect 262916 24080 262922 24132
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 298830 22760 298836 22772
rect 8352 22732 298836 22760
rect 8352 22720 8358 22732
rect 298830 22720 298836 22732
rect 298888 22720 298894 22772
rect 59354 21428 59360 21480
rect 59412 21468 59418 21480
rect 292022 21468 292028 21480
rect 59412 21440 292028 21468
rect 59412 21428 59418 21440
rect 292022 21428 292028 21440
rect 292080 21428 292086 21480
rect 11146 21360 11152 21412
rect 11204 21400 11210 21412
rect 253290 21400 253296 21412
rect 11204 21372 253296 21400
rect 11204 21360 11210 21372
rect 253290 21360 253296 21372
rect 253348 21360 253354 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 32398 20652 32404 20664
rect 3476 20624 32404 20652
rect 3476 20612 3482 20624
rect 32398 20612 32404 20624
rect 32456 20612 32462 20664
rect 216122 20612 216128 20664
rect 216180 20652 216186 20664
rect 579890 20652 579896 20664
rect 216180 20624 579896 20652
rect 216180 20612 216186 20624
rect 579890 20612 579896 20624
rect 579948 20612 579954 20664
rect 175182 20000 175188 20052
rect 175240 20040 175246 20052
rect 262214 20040 262220 20052
rect 175240 20012 262220 20040
rect 175240 20000 175246 20012
rect 262214 20000 262220 20012
rect 262272 20000 262278 20052
rect 91094 19932 91100 19984
rect 91152 19972 91158 19984
rect 283650 19972 283656 19984
rect 91152 19944 283656 19972
rect 91152 19932 91158 19944
rect 283650 19932 283656 19944
rect 283708 19932 283714 19984
rect 114554 18572 114560 18624
rect 114612 18612 114618 18624
rect 283742 18612 283748 18624
rect 114612 18584 283748 18612
rect 114612 18572 114618 18584
rect 283742 18572 283748 18584
rect 283800 18572 283806 18624
rect 187694 17416 187700 17468
rect 187752 17456 187758 17468
rect 253198 17456 253204 17468
rect 187752 17428 253204 17456
rect 187752 17416 187758 17428
rect 253198 17416 253204 17428
rect 253256 17416 253262 17468
rect 207014 17348 207020 17400
rect 207072 17388 207078 17400
rect 345014 17388 345020 17400
rect 207072 17360 345020 17388
rect 207072 17348 207078 17360
rect 345014 17348 345020 17360
rect 345072 17348 345078 17400
rect 95234 17280 95240 17332
rect 95292 17320 95298 17332
rect 302878 17320 302884 17332
rect 95292 17292 302884 17320
rect 95292 17280 95298 17292
rect 302878 17280 302884 17292
rect 302936 17280 302942 17332
rect 24854 17212 24860 17264
rect 24912 17252 24918 17264
rect 256142 17252 256148 17264
rect 24912 17224 256148 17252
rect 24912 17212 24918 17224
rect 256142 17212 256148 17224
rect 256200 17212 256206 17264
rect 112346 15852 112352 15904
rect 112404 15892 112410 15904
rect 305638 15892 305644 15904
rect 112404 15864 305644 15892
rect 112404 15852 112410 15864
rect 305638 15852 305644 15864
rect 305696 15852 305702 15904
rect 179414 14560 179420 14612
rect 179472 14600 179478 14612
rect 306374 14600 306380 14612
rect 179472 14572 306380 14600
rect 179472 14560 179478 14572
rect 306374 14560 306380 14572
rect 306432 14560 306438 14612
rect 122282 14492 122288 14544
rect 122340 14532 122346 14544
rect 256050 14532 256056 14544
rect 122340 14504 256056 14532
rect 122340 14492 122346 14504
rect 256050 14492 256056 14504
rect 256108 14492 256114 14544
rect 66714 14424 66720 14476
rect 66772 14464 66778 14476
rect 293218 14464 293224 14476
rect 66772 14436 293224 14464
rect 66772 14424 66778 14436
rect 293218 14424 293224 14436
rect 293276 14424 293282 14476
rect 119890 13064 119896 13116
rect 119948 13104 119954 13116
rect 264330 13104 264336 13116
rect 119948 13076 264336 13104
rect 119948 13064 119954 13076
rect 264330 13064 264336 13076
rect 264388 13064 264394 13116
rect 179506 11840 179512 11892
rect 179564 11880 179570 11892
rect 294874 11880 294880 11892
rect 179564 11852 294880 11880
rect 179564 11840 179570 11852
rect 294874 11840 294880 11852
rect 294932 11840 294938 11892
rect 109034 11772 109040 11824
rect 109092 11812 109098 11824
rect 265710 11812 265716 11824
rect 109092 11784 265716 11812
rect 109092 11772 109098 11784
rect 265710 11772 265716 11784
rect 265768 11772 265774 11824
rect 33594 11704 33600 11756
rect 33652 11744 33658 11756
rect 292114 11744 292120 11756
rect 33652 11716 292120 11744
rect 33652 11704 33658 11716
rect 292114 11704 292120 11716
rect 292172 11704 292178 11756
rect 106 10956 112 11008
rect 164 10996 170 11008
rect 1302 10996 1308 11008
rect 164 10968 1308 10996
rect 164 10956 170 10968
rect 1302 10956 1308 10968
rect 1360 10996 1366 11008
rect 251174 10996 251180 11008
rect 1360 10968 251180 10996
rect 1360 10956 1366 10968
rect 251174 10956 251180 10968
rect 251232 10956 251238 11008
rect 177942 10344 177948 10396
rect 178000 10384 178006 10396
rect 287330 10384 287336 10396
rect 178000 10356 287336 10384
rect 178000 10344 178006 10356
rect 287330 10344 287336 10356
rect 287388 10344 287394 10396
rect 78122 10276 78128 10328
rect 78180 10316 78186 10328
rect 295978 10316 295984 10328
rect 78180 10288 295984 10316
rect 78180 10276 78186 10288
rect 295978 10276 295984 10288
rect 296036 10276 296042 10328
rect 232498 9052 232504 9104
rect 232556 9092 232562 9104
rect 281902 9092 281908 9104
rect 232556 9064 281908 9092
rect 232556 9052 232562 9064
rect 281902 9052 281908 9064
rect 281960 9052 281966 9104
rect 196618 8984 196624 9036
rect 196676 9024 196682 9036
rect 260650 9024 260656 9036
rect 196676 8996 260656 9024
rect 196676 8984 196682 8996
rect 260650 8984 260656 8996
rect 260708 8984 260714 9036
rect 15930 8916 15936 8968
rect 15988 8956 15994 8968
rect 289078 8956 289084 8968
rect 15988 8928 289084 8956
rect 15988 8916 15994 8928
rect 289078 8916 289084 8928
rect 289136 8916 289142 8968
rect 192478 7692 192484 7744
rect 192536 7732 192542 7744
rect 299658 7732 299664 7744
rect 192536 7704 299664 7732
rect 192536 7692 192542 7704
rect 299658 7692 299664 7704
rect 299716 7692 299722 7744
rect 62022 7624 62028 7676
rect 62080 7664 62086 7676
rect 298738 7664 298744 7676
rect 62080 7636 298744 7664
rect 62080 7624 62086 7636
rect 298738 7624 298744 7636
rect 298796 7624 298802 7676
rect 24210 7556 24216 7608
rect 24268 7596 24274 7608
rect 279418 7596 279424 7608
rect 24268 7568 279424 7596
rect 24268 7556 24274 7568
rect 279418 7556 279424 7568
rect 279476 7556 279482 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 22738 6848 22744 6860
rect 3476 6820 22744 6848
rect 3476 6808 3482 6820
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 260098 6400 260104 6452
rect 260156 6440 260162 6452
rect 284294 6440 284300 6452
rect 260156 6412 284300 6440
rect 260156 6400 260162 6412
rect 284294 6400 284300 6412
rect 284352 6400 284358 6452
rect 206278 6332 206284 6384
rect 206336 6372 206342 6384
rect 266538 6372 266544 6384
rect 206336 6344 266544 6372
rect 206336 6332 206342 6344
rect 266538 6332 266544 6344
rect 266596 6332 266602 6384
rect 198734 6264 198740 6316
rect 198792 6304 198798 6316
rect 276014 6304 276020 6316
rect 198792 6276 276020 6304
rect 198792 6264 198798 6276
rect 276014 6264 276020 6276
rect 276072 6264 276078 6316
rect 31662 6196 31668 6248
rect 31720 6236 31726 6248
rect 136450 6236 136456 6248
rect 31720 6208 136456 6236
rect 31720 6196 31726 6208
rect 136450 6196 136456 6208
rect 136508 6196 136514 6248
rect 197998 6196 198004 6248
rect 198056 6236 198062 6248
rect 292574 6236 292580 6248
rect 198056 6208 292580 6236
rect 198056 6196 198062 6208
rect 292574 6196 292580 6208
rect 292632 6196 292638 6248
rect 70302 6128 70308 6180
rect 70360 6168 70366 6180
rect 301498 6168 301504 6180
rect 70360 6140 301504 6168
rect 70360 6128 70366 6140
rect 301498 6128 301504 6140
rect 301556 6128 301562 6180
rect 305546 6128 305552 6180
rect 305604 6168 305610 6180
rect 338114 6168 338120 6180
rect 305604 6140 338120 6168
rect 305604 6128 305610 6140
rect 338114 6128 338120 6140
rect 338172 6128 338178 6180
rect 193214 4904 193220 4956
rect 193272 4944 193278 4956
rect 247586 4944 247592 4956
rect 193272 4916 247592 4944
rect 193272 4904 193278 4916
rect 247586 4904 247592 4916
rect 247644 4904 247650 4956
rect 249978 4904 249984 4956
rect 250036 4944 250042 4956
rect 265618 4944 265624 4956
rect 250036 4916 265624 4944
rect 250036 4904 250042 4916
rect 265618 4904 265624 4916
rect 265676 4904 265682 4956
rect 175090 4836 175096 4888
rect 175148 4876 175154 4888
rect 304350 4876 304356 4888
rect 175148 4848 304356 4876
rect 175148 4836 175154 4848
rect 304350 4836 304356 4848
rect 304408 4836 304414 4888
rect 48958 4768 48964 4820
rect 49016 4808 49022 4820
rect 278130 4808 278136 4820
rect 49016 4780 278136 4808
rect 49016 4768 49022 4780
rect 278130 4768 278136 4780
rect 278188 4768 278194 4820
rect 335998 4156 336004 4208
rect 336056 4196 336062 4208
rect 340966 4196 340972 4208
rect 336056 4168 340972 4196
rect 336056 4156 336062 4168
rect 340966 4156 340972 4168
rect 341024 4156 341030 4208
rect 261570 4088 261576 4140
rect 261628 4128 261634 4140
rect 268838 4128 268844 4140
rect 261628 4100 268844 4128
rect 261628 4088 261634 4100
rect 268838 4088 268844 4100
rect 268896 4088 268902 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 316218 4128 316224 4140
rect 315356 4100 316224 4128
rect 315356 4088 315362 4100
rect 316218 4088 316224 4100
rect 316276 4088 316282 4140
rect 211798 3748 211804 3800
rect 211856 3788 211862 3800
rect 245194 3788 245200 3800
rect 211856 3760 245200 3788
rect 211856 3748 211862 3760
rect 245194 3748 245200 3760
rect 245252 3748 245258 3800
rect 204898 3680 204904 3732
rect 204956 3720 204962 3732
rect 242894 3720 242900 3732
rect 204956 3692 242900 3720
rect 204956 3680 204962 3692
rect 242894 3680 242900 3692
rect 242952 3680 242958 3732
rect 264882 3680 264888 3732
rect 264940 3720 264946 3732
rect 271230 3720 271236 3732
rect 264940 3692 271236 3720
rect 264940 3680 264946 3692
rect 271230 3680 271236 3692
rect 271288 3680 271294 3732
rect 204162 3612 204168 3664
rect 204220 3652 204226 3664
rect 248782 3652 248788 3664
rect 204220 3624 248788 3652
rect 204220 3612 204226 3624
rect 248782 3612 248788 3624
rect 248840 3612 248846 3664
rect 253198 3612 253204 3664
rect 253256 3652 253262 3664
rect 261754 3652 261760 3664
rect 253256 3624 261760 3652
rect 253256 3612 253262 3624
rect 261754 3612 261760 3624
rect 261812 3612 261818 3664
rect 268378 3612 268384 3664
rect 268436 3652 268442 3664
rect 283098 3652 283104 3664
rect 268436 3624 283104 3652
rect 268436 3612 268442 3624
rect 283098 3612 283104 3624
rect 283156 3612 283162 3664
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 56594 3584 56600 3596
rect 6512 3556 56600 3584
rect 6512 3544 6518 3556
rect 56594 3544 56600 3556
rect 56652 3544 56658 3596
rect 102134 3544 102140 3596
rect 102192 3584 102198 3596
rect 103330 3584 103336 3596
rect 102192 3556 103336 3584
rect 102192 3544 102198 3556
rect 103330 3544 103336 3556
rect 103388 3544 103394 3596
rect 123478 3544 123484 3596
rect 123536 3584 123542 3596
rect 228358 3584 228364 3596
rect 123536 3556 228364 3584
rect 123536 3544 123542 3556
rect 228358 3544 228364 3556
rect 228416 3544 228422 3596
rect 244090 3544 244096 3596
rect 244148 3584 244154 3596
rect 255958 3584 255964 3596
rect 244148 3556 255964 3584
rect 244148 3544 244154 3556
rect 255958 3544 255964 3556
rect 256016 3544 256022 3596
rect 259454 3544 259460 3596
rect 259512 3584 259518 3596
rect 275278 3584 275284 3596
rect 259512 3556 275284 3584
rect 259512 3544 259518 3556
rect 275278 3544 275284 3556
rect 275336 3544 275342 3596
rect 278038 3544 278044 3596
rect 278096 3584 278102 3596
rect 288986 3584 288992 3596
rect 278096 3556 288992 3584
rect 278096 3544 278102 3556
rect 288986 3544 288992 3556
rect 289044 3544 289050 3596
rect 289722 3544 289728 3596
rect 289780 3584 289786 3596
rect 293678 3584 293684 3596
rect 289780 3556 293684 3584
rect 289780 3544 289786 3556
rect 293678 3544 293684 3556
rect 293736 3544 293742 3596
rect 323578 3544 323584 3596
rect 323636 3584 323642 3596
rect 337470 3584 337476 3596
rect 323636 3556 337476 3584
rect 323636 3544 323642 3556
rect 337470 3544 337476 3556
rect 337528 3544 337534 3596
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 20254 3516 20260 3528
rect 19392 3488 20260 3516
rect 19392 3476 19398 3488
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36814 3516 36820 3528
rect 35952 3488 36820 3516
rect 35952 3476 35958 3488
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53374 3516 53380 3528
rect 52512 3488 53380 3516
rect 52512 3476 52518 3488
rect 53374 3476 53380 3488
rect 53432 3476 53438 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 185578 3516 185584 3528
rect 57296 3488 185584 3516
rect 57296 3476 57302 3488
rect 185578 3476 185584 3488
rect 185636 3476 185642 3528
rect 189718 3476 189724 3528
rect 189776 3516 189782 3528
rect 240502 3516 240508 3528
rect 189776 3488 240508 3516
rect 189776 3476 189782 3488
rect 240502 3476 240508 3488
rect 240560 3476 240566 3528
rect 252370 3476 252376 3528
rect 252428 3516 252434 3528
rect 270494 3516 270500 3528
rect 252428 3488 270500 3516
rect 252428 3476 252434 3488
rect 270494 3476 270500 3488
rect 270552 3476 270558 3528
rect 280798 3516 280804 3528
rect 277366 3488 280804 3516
rect 28902 3408 28908 3460
rect 28960 3448 28966 3460
rect 214558 3448 214564 3460
rect 28960 3420 214564 3448
rect 28960 3408 28966 3420
rect 214558 3408 214564 3420
rect 214616 3408 214622 3460
rect 215938 3408 215944 3460
rect 215996 3448 216002 3460
rect 254670 3448 254676 3460
rect 215996 3420 254676 3448
rect 215996 3408 216002 3420
rect 254670 3408 254676 3420
rect 254728 3408 254734 3460
rect 264146 3408 264152 3460
rect 264204 3448 264210 3460
rect 277366 3448 277394 3488
rect 280798 3476 280804 3488
rect 280856 3476 280862 3528
rect 287698 3476 287704 3528
rect 287756 3516 287762 3528
rect 291378 3516 291384 3528
rect 287756 3488 291384 3516
rect 287756 3476 287762 3488
rect 291378 3476 291384 3488
rect 291436 3476 291442 3528
rect 299474 3476 299480 3528
rect 299532 3516 299538 3528
rect 300762 3516 300768 3528
rect 299532 3488 300768 3516
rect 299532 3476 299538 3488
rect 300762 3476 300768 3488
rect 300820 3476 300826 3528
rect 316126 3476 316132 3528
rect 316184 3516 316190 3528
rect 317322 3516 317328 3528
rect 316184 3488 317328 3516
rect 316184 3476 316190 3488
rect 317322 3476 317328 3488
rect 317380 3476 317386 3528
rect 324406 3476 324412 3528
rect 324464 3516 324470 3528
rect 325602 3516 325608 3528
rect 324464 3488 325608 3516
rect 324464 3476 324470 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 332594 3476 332600 3528
rect 332652 3516 332658 3528
rect 333882 3516 333888 3528
rect 332652 3488 333888 3516
rect 332652 3476 332658 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 340874 3516 340880 3528
rect 334084 3488 340880 3516
rect 264204 3420 277394 3448
rect 264204 3408 264210 3420
rect 280706 3408 280712 3460
rect 280764 3448 280770 3460
rect 282178 3448 282184 3460
rect 280764 3420 282184 3448
rect 280764 3408 280770 3420
rect 282178 3408 282184 3420
rect 282236 3408 282242 3460
rect 291838 3408 291844 3460
rect 291896 3448 291902 3460
rect 298462 3448 298468 3460
rect 291896 3420 298468 3448
rect 291896 3408 291902 3420
rect 298462 3408 298468 3420
rect 298520 3408 298526 3460
rect 309778 3408 309784 3460
rect 309836 3448 309842 3460
rect 322106 3448 322112 3460
rect 309836 3420 322112 3448
rect 309836 3408 309842 3420
rect 322106 3408 322112 3420
rect 322164 3408 322170 3460
rect 326798 3340 326804 3392
rect 326856 3380 326862 3392
rect 334084 3380 334112 3488
rect 340874 3476 340880 3488
rect 340932 3476 340938 3528
rect 326856 3352 334112 3380
rect 326856 3340 326862 3352
rect 323302 3272 323308 3324
rect 323360 3312 323366 3324
rect 342254 3312 342260 3324
rect 323360 3284 342260 3312
rect 323360 3272 323366 3284
rect 342254 3272 342260 3284
rect 342312 3272 342318 3324
rect 264238 3204 264244 3256
rect 264296 3244 264302 3256
rect 270034 3244 270040 3256
rect 264296 3216 270040 3244
rect 264296 3204 264302 3216
rect 270034 3204 270040 3216
rect 270092 3204 270098 3256
rect 330386 3204 330392 3256
rect 330444 3244 330450 3256
rect 331490 3244 331496 3256
rect 330444 3216 331496 3244
rect 330444 3204 330450 3216
rect 331490 3204 331496 3216
rect 331548 3204 331554 3256
rect 308490 3136 308496 3188
rect 308548 3176 308554 3188
rect 315022 3176 315028 3188
rect 308548 3148 315028 3176
rect 308548 3136 308554 3148
rect 315022 3136 315028 3148
rect 315080 3136 315086 3188
rect 345658 3136 345664 3188
rect 345716 3176 345722 3188
rect 349246 3176 349252 3188
rect 345716 3148 349252 3176
rect 345716 3136 345722 3148
rect 349246 3136 349252 3148
rect 349304 3136 349310 3188
rect 249702 3000 249708 3052
rect 249760 3040 249766 3052
rect 255866 3040 255872 3052
rect 249760 3012 255872 3040
rect 249760 3000 249766 3012
rect 255866 3000 255872 3012
rect 255924 3000 255930 3052
rect 235810 2932 235816 2984
rect 235868 2972 235874 2984
rect 238018 2972 238024 2984
rect 235868 2944 238024 2972
rect 235868 2932 235874 2944
rect 238018 2932 238024 2944
rect 238076 2932 238082 2984
rect 337378 2932 337384 2984
rect 337436 2972 337442 2984
rect 338666 2972 338672 2984
rect 337436 2944 338672 2972
rect 337436 2932 337442 2944
rect 338666 2932 338672 2944
rect 338724 2932 338730 2984
rect 56042 2048 56048 2100
rect 56100 2088 56106 2100
rect 297450 2088 297456 2100
rect 56100 2060 297456 2088
rect 56100 2048 56106 2060
rect 297450 2048 297456 2060
rect 297508 2048 297514 2100
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 37188 702788 37240 702840
rect 202788 702788 202840 702840
rect 63408 702720 63460 702772
rect 267648 702720 267700 702772
rect 297364 702720 297416 702772
rect 494796 702720 494848 702772
rect 8116 702652 8168 702704
rect 210424 702652 210476 702704
rect 248328 702652 248380 702704
rect 527180 702652 527232 702704
rect 130384 702584 130436 702636
rect 413652 702584 413704 702636
rect 53748 702516 53800 702568
rect 462320 702516 462372 702568
rect 63316 702448 63368 702500
rect 543464 702448 543516 702500
rect 24308 700340 24360 700392
rect 48964 700340 49016 700392
rect 45468 700272 45520 700324
rect 137836 700272 137888 700324
rect 235172 700272 235224 700324
rect 244280 700272 244332 700324
rect 253204 700272 253256 700324
rect 559656 700272 559708 700324
rect 100024 699660 100076 699712
rect 105452 699660 105504 699712
rect 395344 699660 395396 699712
rect 397460 699660 397512 699712
rect 63500 698912 63552 698964
rect 218980 698912 219032 698964
rect 262128 698912 262180 698964
rect 429844 698912 429896 698964
rect 278044 697552 278096 697604
rect 348792 697552 348844 697604
rect 363604 696940 363656 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 46204 683136 46256 683188
rect 242808 683136 242860 683188
rect 580172 683136 580224 683188
rect 291844 670692 291896 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 43444 656888 43496 656940
rect 251088 643084 251140 643136
rect 580172 643084 580224 643136
rect 3516 632068 3568 632120
rect 229744 632068 229796 632120
rect 175372 630640 175424 630692
rect 244372 630640 244424 630692
rect 580172 630640 580224 630692
rect 3516 618604 3568 618656
rect 7564 618604 7616 618656
rect 48964 607112 49016 607164
rect 52276 607112 52328 607164
rect 3516 606024 3568 606076
rect 8944 606024 8996 606076
rect 52276 605820 52328 605872
rect 185032 605820 185084 605872
rect 88340 600924 88392 600976
rect 236644 600924 236696 600976
rect 71780 599564 71832 599616
rect 245752 599564 245804 599616
rect 40040 596776 40092 596828
rect 217324 596776 217376 596828
rect 169760 595416 169812 595468
rect 245844 595416 245896 595468
rect 3424 594056 3476 594108
rect 244556 594056 244608 594108
rect 256608 594056 256660 594108
rect 299480 594056 299532 594108
rect 90180 592628 90232 592680
rect 100024 592628 100076 592680
rect 220728 592628 220780 592680
rect 282920 592628 282972 592680
rect 46848 592152 46900 592204
rect 102600 592152 102652 592204
rect 45284 592084 45336 592136
rect 134156 592084 134208 592136
rect 48136 592016 48188 592068
rect 153476 592016 153528 592068
rect 153200 591268 153252 591320
rect 251180 591268 251232 591320
rect 53656 590860 53708 590912
rect 86500 590860 86552 590912
rect 42616 590792 42668 590844
rect 112260 590792 112312 590844
rect 44088 590724 44140 590776
rect 143816 590724 143868 590776
rect 46756 590656 46808 590708
rect 159916 590656 159968 590708
rect 130384 590248 130436 590300
rect 130936 590248 130988 590300
rect 201408 589908 201460 589960
rect 580172 589908 580224 589960
rect 55036 589636 55088 589688
rect 118700 589636 118752 589688
rect 53564 589568 53616 589620
rect 121920 589568 121972 589620
rect 61936 589500 61988 589552
rect 130936 589500 130988 589552
rect 52184 589432 52236 589484
rect 140596 589432 140648 589484
rect 42708 589364 42760 589416
rect 156696 589364 156748 589416
rect 35808 589296 35860 589348
rect 163136 589296 163188 589348
rect 236000 589296 236052 589348
rect 236644 589296 236696 589348
rect 258080 589296 258132 589348
rect 256700 588548 256752 588600
rect 331220 588548 331272 588600
rect 56416 588208 56468 588260
rect 90180 588208 90232 588260
rect 39672 588140 39724 588192
rect 105912 588140 105964 588192
rect 229744 588140 229796 588192
rect 249800 588140 249852 588192
rect 60096 588072 60148 588124
rect 127808 588072 127860 588124
rect 226340 588072 226392 588124
rect 256700 588072 256752 588124
rect 54944 588004 54996 588056
rect 191564 588004 191616 588056
rect 210424 588004 210476 588056
rect 244464 588004 244516 588056
rect 5448 587936 5500 587988
rect 147128 587936 147180 587988
rect 242808 587936 242860 587988
rect 289084 587936 289136 587988
rect 48964 587868 49016 587920
rect 198004 587868 198056 587920
rect 246304 587868 246356 587920
rect 35164 586916 35216 586968
rect 80152 586916 80204 586968
rect 34428 586848 34480 586900
rect 77576 586848 77628 586900
rect 239220 586848 239272 586900
rect 252560 586848 252612 586900
rect 49516 586780 49568 586832
rect 96252 586780 96304 586832
rect 217324 586780 217376 586832
rect 243176 586780 243228 586832
rect 60004 586712 60056 586764
rect 109132 586712 109184 586764
rect 214104 586712 214156 586764
rect 248420 586712 248472 586764
rect 62764 586644 62816 586696
rect 115572 586644 115624 586696
rect 207664 586644 207716 586696
rect 255320 586644 255372 586696
rect 79416 586576 79468 586628
rect 137468 586576 137520 586628
rect 181904 586576 181956 586628
rect 242992 586576 243044 586628
rect 63592 586508 63644 586560
rect 150348 586508 150400 586560
rect 172888 586508 172940 586560
rect 259460 586508 259512 586560
rect 63224 585760 63276 585812
rect 79416 585760 79468 585812
rect 44824 585420 44876 585472
rect 71136 585420 71188 585472
rect 41236 585352 41288 585404
rect 67916 585352 67968 585404
rect 194784 585352 194836 585404
rect 243636 585352 243688 585404
rect 251916 585352 251968 585404
rect 50344 585284 50396 585336
rect 172888 585284 172940 585336
rect 220544 585284 220596 585336
rect 220728 585284 220780 585336
rect 292580 585284 292632 585336
rect 31024 585216 31076 585268
rect 263692 585216 263744 585268
rect 52368 585148 52420 585200
rect 125232 585148 125284 585200
rect 166448 585148 166500 585200
rect 245660 585148 245712 585200
rect 57888 583856 57940 583908
rect 63592 583856 63644 583908
rect 49608 583788 49660 583840
rect 73988 584536 74040 584588
rect 204720 584536 204772 584588
rect 251272 583788 251324 583840
rect 2872 583720 2924 583772
rect 57704 583720 57756 583772
rect 57888 583720 57940 583772
rect 58716 583720 58768 583772
rect 247132 583720 247184 583772
rect 245660 582360 245712 582412
rect 336740 582360 336792 582412
rect 243176 581612 243228 581664
rect 276020 581612 276072 581664
rect 243268 578144 243320 578196
rect 579804 578144 579856 578196
rect 245752 576512 245804 576564
rect 245936 576512 245988 576564
rect 245752 575492 245804 575544
rect 335360 575492 335412 575544
rect 245752 572704 245804 572756
rect 287704 572704 287756 572756
rect 55128 568556 55180 568608
rect 60740 568556 60792 568608
rect 3424 565836 3476 565888
rect 14464 565836 14516 565888
rect 245752 565836 245804 565888
rect 332600 565836 332652 565888
rect 27528 564408 27580 564460
rect 60740 564408 60792 564460
rect 445024 563048 445076 563100
rect 580172 563048 580224 563100
rect 48228 561688 48280 561740
rect 60740 561688 60792 561740
rect 245752 558900 245804 558952
rect 248512 558900 248564 558952
rect 245752 556180 245804 556232
rect 314660 556180 314712 556232
rect 500224 556180 500276 556232
rect 33048 554752 33100 554804
rect 60740 554752 60792 554804
rect 3148 554684 3200 554736
rect 31024 554684 31076 554736
rect 39856 552032 39908 552084
rect 60740 552032 60792 552084
rect 264980 549856 265032 549908
rect 363604 549856 363656 549908
rect 245752 549244 245804 549296
rect 264980 549244 265032 549296
rect 57888 548360 57940 548412
rect 60740 548360 60792 548412
rect 7564 542988 7616 543040
rect 39948 542988 40000 543040
rect 39948 542376 40000 542428
rect 60740 542376 60792 542428
rect 245752 539588 245804 539640
rect 328460 539588 328512 539640
rect 245752 539452 245804 539504
rect 245936 539452 245988 539504
rect 31576 538228 31628 538280
rect 60740 538228 60792 538280
rect 257344 536800 257396 536852
rect 579896 536800 579948 536852
rect 245844 536052 245896 536104
rect 313280 536052 313332 536104
rect 57244 535440 57296 535492
rect 60740 535440 60792 535492
rect 242992 532720 243044 532772
rect 243268 532720 243320 532772
rect 46204 529864 46256 529916
rect 53472 529864 53524 529916
rect 53472 528572 53524 528624
rect 60740 528572 60792 528624
rect 3700 527144 3752 527196
rect 4068 527144 4120 527196
rect 46204 527144 46256 527196
rect 245844 525784 245896 525836
rect 282184 525784 282236 525836
rect 59176 521636 59228 521688
rect 61660 521636 61712 521688
rect 245844 521636 245896 521688
rect 349252 521636 349304 521688
rect 245844 518916 245896 518968
rect 259552 518916 259604 518968
rect 3424 516060 3476 516112
rect 58716 516060 58768 516112
rect 38568 514768 38620 514820
rect 60740 514768 60792 514820
rect 245384 514768 245436 514820
rect 263600 514768 263652 514820
rect 58716 513884 58768 513936
rect 60096 513884 60148 513936
rect 245844 512592 245896 512644
rect 251088 512592 251140 512644
rect 296720 512592 296772 512644
rect 251824 510620 251876 510672
rect 580172 510620 580224 510672
rect 246672 509804 246724 509856
rect 248328 509804 248380 509856
rect 248328 509260 248380 509312
rect 249892 509260 249944 509312
rect 245844 506404 245896 506456
rect 263692 506404 263744 506456
rect 263692 505724 263744 505776
rect 300860 505724 300912 505776
rect 245844 502324 245896 502376
rect 324964 502324 325016 502376
rect 3056 500964 3108 501016
rect 50436 500964 50488 501016
rect 55864 500964 55916 501016
rect 60740 500964 60792 501016
rect 245844 499536 245896 499588
rect 329840 499536 329892 499588
rect 262128 496816 262180 496868
rect 305000 496816 305052 496868
rect 245844 496748 245896 496800
rect 48044 495456 48096 495508
rect 60740 495456 60792 495508
rect 245844 492668 245896 492720
rect 270500 492668 270552 492720
rect 56232 491308 56284 491360
rect 60740 491308 60792 491360
rect 32956 488520 33008 488572
rect 60740 488520 60792 488572
rect 43996 485800 44048 485852
rect 61200 485800 61252 485852
rect 245844 485800 245896 485852
rect 261484 485800 261536 485852
rect 251916 485732 251968 485784
rect 580172 485732 580224 485784
rect 251088 482264 251140 482316
rect 580264 482264 580316 482316
rect 59084 481652 59136 481704
rect 61568 481652 61620 481704
rect 13084 477504 13136 477556
rect 60740 477504 60792 477556
rect 3424 474716 3476 474768
rect 22744 474716 22796 474768
rect 245844 474716 245896 474768
rect 317420 474716 317472 474768
rect 299480 472608 299532 472660
rect 364340 472608 364392 472660
rect 245844 471996 245896 472048
rect 299480 471996 299532 472048
rect 45376 470568 45428 470620
rect 60924 470568 60976 470620
rect 275284 470568 275336 470620
rect 580080 470568 580132 470620
rect 37096 467848 37148 467900
rect 60740 467848 60792 467900
rect 53748 464992 53800 465044
rect 60740 464992 60792 465044
rect 3424 463632 3476 463684
rect 50344 463632 50396 463684
rect 17224 460912 17276 460964
rect 52092 460912 52144 460964
rect 60740 460912 60792 460964
rect 245936 460912 245988 460964
rect 269764 460912 269816 460964
rect 245936 458804 245988 458856
rect 249984 458804 250036 458856
rect 50804 456764 50856 456816
rect 60740 456764 60792 456816
rect 249064 456764 249116 456816
rect 580172 456764 580224 456816
rect 245936 455404 245988 455456
rect 263692 455404 263744 455456
rect 60648 455336 60700 455388
rect 61384 455336 61436 455388
rect 246304 450508 246356 450560
rect 252652 450508 252704 450560
rect 63224 449896 63276 449948
rect 63500 449896 63552 449948
rect 3332 449828 3384 449880
rect 17224 449828 17276 449880
rect 245936 448536 245988 448588
rect 255412 448536 255464 448588
rect 245384 447040 245436 447092
rect 278044 447040 278096 447092
rect 54852 444388 54904 444440
rect 60740 444388 60792 444440
rect 50896 441600 50948 441652
rect 60740 441600 60792 441652
rect 245936 438880 245988 438932
rect 278044 438880 278096 438932
rect 46664 437452 46716 437504
rect 60924 437452 60976 437504
rect 59268 434732 59320 434784
rect 61568 434732 61620 434784
rect 245936 434732 245988 434784
rect 327264 434732 327316 434784
rect 57704 433236 57756 433288
rect 62856 433236 62908 433288
rect 245936 433236 245988 433288
rect 251088 433304 251140 433356
rect 306380 433304 306432 433356
rect 22744 428408 22796 428460
rect 49424 428408 49476 428460
rect 49424 427796 49476 427848
rect 60740 427796 60792 427848
rect 245936 427796 245988 427848
rect 291936 427796 291988 427848
rect 252468 425688 252520 425740
rect 291844 425688 291896 425740
rect 245936 425076 245988 425128
rect 251364 425076 251416 425128
rect 252468 425076 252520 425128
rect 39764 423648 39816 423700
rect 60740 423648 60792 423700
rect 245936 420928 245988 420980
rect 322940 420928 322992 420980
rect 500224 419432 500276 419484
rect 580172 419432 580224 419484
rect 245936 418208 245988 418260
rect 247316 418208 247368 418260
rect 58992 417392 59044 417444
rect 60004 417392 60056 417444
rect 62856 417392 62908 417444
rect 63132 417392 63184 417444
rect 17224 416780 17276 416832
rect 62304 416780 62356 416832
rect 63224 416780 63276 416832
rect 60464 416712 60516 416764
rect 62764 416712 62816 416764
rect 42524 413992 42576 414044
rect 60740 413992 60792 414044
rect 245936 413992 245988 414044
rect 292764 413992 292816 414044
rect 245936 411272 245988 411324
rect 298192 411272 298244 411324
rect 3424 411204 3476 411256
rect 48964 411204 49016 411256
rect 53564 409980 53616 410032
rect 53748 409980 53800 410032
rect 245292 408484 245344 408536
rect 310612 408484 310664 408536
rect 37188 407736 37240 407788
rect 60740 407736 60792 407788
rect 249156 407736 249208 407788
rect 580356 407736 580408 407788
rect 243084 407124 243136 407176
rect 245660 407124 245712 407176
rect 3516 407056 3568 407108
rect 7840 407056 7892 407108
rect 7840 405696 7892 405748
rect 8208 405696 8260 405748
rect 57336 405696 57388 405748
rect 53748 405084 53800 405136
rect 66904 405084 66956 405136
rect 236644 405084 236696 405136
rect 260840 405084 260892 405136
rect 56416 405016 56468 405068
rect 80060 405016 80112 405068
rect 171048 405016 171100 405068
rect 243084 405016 243136 405068
rect 57704 404948 57756 405000
rect 104164 404948 104216 405000
rect 165528 404948 165580 405000
rect 249892 404948 249944 405000
rect 8944 404472 8996 404524
rect 96528 404472 96580 404524
rect 120724 404472 120776 404524
rect 202880 404472 202932 404524
rect 203800 404472 203852 404524
rect 251824 404472 251876 404524
rect 50436 404404 50488 404456
rect 178040 404404 178092 404456
rect 197360 404404 197412 404456
rect 249064 404404 249116 404456
rect 66168 404336 66220 404388
rect 580172 404336 580224 404388
rect 105268 404268 105320 404320
rect 445024 404268 445076 404320
rect 14464 404200 14516 404252
rect 242164 404200 242216 404252
rect 222844 404132 222896 404184
rect 257344 404132 257396 404184
rect 63500 403996 63552 404048
rect 63960 403996 64012 404048
rect 50988 403792 51040 403844
rect 68284 403792 68336 403844
rect 55036 403724 55088 403776
rect 73804 403724 73856 403776
rect 60372 403656 60424 403708
rect 98736 403656 98788 403708
rect 239404 403656 239456 403708
rect 248420 403656 248472 403708
rect 63132 403588 63184 403640
rect 124220 403588 124272 403640
rect 148416 403588 148468 403640
rect 251272 403588 251324 403640
rect 240140 403520 240192 403572
rect 244464 403520 244516 403572
rect 46204 402908 46256 402960
rect 200764 402908 200816 402960
rect 209596 402908 209648 402960
rect 256608 402908 256660 402960
rect 57336 402840 57388 402892
rect 181444 402840 181496 402892
rect 43444 402772 43496 402824
rect 79324 402772 79376 402824
rect 161940 402772 161992 402824
rect 162768 402772 162820 402824
rect 249156 402772 249208 402824
rect 100668 402296 100720 402348
rect 108488 402296 108540 402348
rect 117504 402296 117556 402348
rect 126980 402296 127032 402348
rect 164148 402296 164200 402348
rect 171600 402296 171652 402348
rect 193864 402296 193916 402348
rect 252652 402296 252704 402348
rect 256608 402296 256660 402348
rect 299572 402296 299624 402348
rect 102048 402228 102100 402280
rect 122104 402228 122156 402280
rect 136824 402228 136876 402280
rect 146300 402228 146352 402280
rect 168288 402228 168340 402280
rect 197360 402228 197412 402280
rect 232136 402228 232188 402280
rect 309140 402228 309192 402280
rect 102784 401752 102836 401804
rect 105268 401752 105320 401804
rect 116584 401616 116636 401668
rect 123944 401616 123996 401668
rect 127164 401616 127216 401668
rect 129004 401616 129056 401668
rect 158076 401616 158128 401668
rect 158720 401616 158772 401668
rect 214564 401004 214616 401056
rect 247316 401004 247368 401056
rect 177856 400936 177908 400988
rect 242992 400936 243044 400988
rect 48136 400868 48188 400920
rect 82084 400868 82136 400920
rect 173716 400868 173768 400920
rect 255320 400868 255372 400920
rect 82728 400120 82780 400172
rect 477500 400120 477552 400172
rect 53564 400052 53616 400104
rect 296812 400052 296864 400104
rect 297364 400052 297416 400104
rect 173808 399576 173860 399628
rect 187700 399576 187752 399628
rect 52276 399508 52328 399560
rect 84844 399508 84896 399560
rect 111064 399508 111116 399560
rect 136640 399508 136692 399560
rect 156604 399508 156656 399560
rect 174820 399508 174872 399560
rect 179788 399508 179840 399560
rect 206376 399508 206428 399560
rect 61752 399440 61804 399492
rect 120724 399440 120776 399492
rect 145564 399440 145616 399492
rect 259552 399440 259604 399492
rect 95148 398760 95200 398812
rect 96528 398760 96580 398812
rect 123484 398148 123536 398200
rect 194140 398148 194192 398200
rect 194600 398148 194652 398200
rect 256700 398148 256752 398200
rect 3976 398080 4028 398132
rect 5448 398080 5500 398132
rect 25504 398080 25556 398132
rect 170956 398080 171008 398132
rect 251364 398080 251416 398132
rect 39672 396924 39724 396976
rect 64144 396924 64196 396976
rect 135904 396924 135956 396976
rect 168380 396924 168432 396976
rect 45284 396856 45336 396908
rect 75184 396856 75236 396908
rect 153108 396856 153160 396908
rect 190920 396856 190972 396908
rect 63224 396788 63276 396840
rect 98644 396788 98696 396840
rect 157984 396788 158036 396840
rect 240140 396788 240192 396840
rect 59084 396720 59136 396772
rect 140780 396720 140832 396772
rect 582380 396720 582432 396772
rect 202144 395428 202196 395480
rect 247224 395428 247276 395480
rect 175188 395360 175240 395412
rect 249800 395360 249852 395412
rect 52184 395292 52236 395344
rect 86224 395292 86276 395344
rect 148324 395292 148376 395344
rect 245844 395292 245896 395344
rect 319444 395292 319496 395344
rect 45284 394000 45336 394052
rect 85580 394000 85632 394052
rect 181444 394000 181496 394052
rect 241520 394000 241572 394052
rect 48136 393932 48188 393984
rect 95240 393932 95292 393984
rect 124864 393932 124916 393984
rect 224960 393932 225012 393984
rect 246304 393320 246356 393372
rect 315304 393320 315356 393372
rect 166264 392640 166316 392692
rect 246304 392640 246356 392692
rect 176476 392572 176528 392624
rect 258080 392572 258132 392624
rect 149704 391960 149756 392012
rect 212540 391960 212592 392012
rect 246396 391960 246448 392012
rect 353300 391960 353352 392012
rect 44088 391280 44140 391332
rect 88340 391280 88392 391332
rect 212540 391280 212592 391332
rect 256700 391280 256752 391332
rect 52368 391212 52420 391264
rect 98000 391212 98052 391264
rect 153844 391212 153896 391264
rect 246396 391212 246448 391264
rect 41144 388424 41196 388476
rect 75920 388424 75972 388476
rect 178040 388288 178092 388340
rect 178684 388288 178736 388340
rect 162124 388220 162176 388272
rect 162768 388220 162820 388272
rect 135996 387880 136048 387932
rect 178040 387880 178092 387932
rect 162768 387812 162820 387864
rect 293960 387812 294012 387864
rect 45468 387744 45520 387796
rect 113180 387744 113232 387796
rect 114468 387744 114520 387796
rect 114468 387064 114520 387116
rect 293040 387064 293092 387116
rect 234620 385636 234672 385688
rect 323032 385636 323084 385688
rect 242164 384344 242216 384396
rect 262220 384344 262272 384396
rect 79324 384276 79376 384328
rect 121460 384276 121512 384328
rect 132408 384276 132460 384328
rect 245752 384276 245804 384328
rect 121460 383664 121512 383716
rect 234620 383664 234672 383716
rect 63868 382916 63920 382968
rect 138020 382916 138072 382968
rect 138020 382236 138072 382288
rect 273904 382236 273956 382288
rect 275284 382236 275336 382288
rect 178684 381556 178736 381608
rect 294052 381556 294104 381608
rect 126244 381488 126296 381540
rect 255412 381488 255464 381540
rect 271328 379448 271380 379500
rect 580172 379448 580224 379500
rect 217324 378768 217376 378820
rect 270500 378768 270552 378820
rect 271328 378768 271380 378820
rect 218060 378088 218112 378140
rect 251180 378088 251232 378140
rect 252468 378088 252520 378140
rect 60556 377408 60608 377460
rect 109684 377408 109736 377460
rect 166816 377408 166868 377460
rect 248512 377408 248564 377460
rect 252468 377408 252520 377460
rect 270500 377408 270552 377460
rect 278044 377408 278096 377460
rect 287060 377408 287112 377460
rect 220084 376048 220136 376100
rect 247040 376048 247092 376100
rect 111708 375980 111760 376032
rect 236644 375980 236696 376032
rect 91100 375300 91152 375352
rect 92388 375300 92440 375352
rect 160836 374620 160888 374672
rect 264980 374620 265032 374672
rect 92388 374008 92440 374060
rect 295616 374008 295668 374060
rect 205640 373328 205692 373380
rect 253204 373328 253256 373380
rect 59176 373260 59228 373312
rect 113824 373260 113876 373312
rect 137284 373260 137336 373312
rect 183560 373260 183612 373312
rect 231124 373260 231176 373312
rect 261484 373260 261536 373312
rect 295524 373260 295576 373312
rect 164240 372580 164292 372632
rect 164884 372580 164936 372632
rect 356060 372580 356112 372632
rect 43904 372172 43956 372224
rect 44824 372172 44876 372224
rect 53656 371900 53708 371952
rect 112444 371900 112496 371952
rect 209044 371900 209096 371952
rect 217324 371900 217376 371952
rect 49424 371832 49476 371884
rect 129832 371832 129884 371884
rect 215300 371832 215352 371884
rect 279424 371832 279476 371884
rect 282184 371832 282236 371884
rect 295340 371832 295392 371884
rect 3424 371220 3476 371272
rect 43904 371220 43956 371272
rect 129832 371220 129884 371272
rect 202972 371220 203024 371272
rect 200764 370608 200816 370660
rect 264980 370608 265032 370660
rect 168196 370540 168248 370592
rect 239404 370540 239456 370592
rect 139308 370472 139360 370524
rect 227720 370472 227772 370524
rect 243360 369180 243412 369232
rect 252560 369180 252612 369232
rect 178684 369112 178736 369164
rect 237380 369112 237432 369164
rect 294144 369112 294196 369164
rect 39672 368500 39724 368552
rect 242992 368500 243044 368552
rect 243360 368500 243412 368552
rect 211804 367820 211856 367872
rect 244556 367820 244608 367872
rect 129740 367752 129792 367804
rect 143540 367752 143592 367804
rect 144276 367752 144328 367804
rect 169116 367752 169168 367804
rect 263692 367752 263744 367804
rect 144276 367072 144328 367124
rect 205640 367072 205692 367124
rect 52092 366392 52144 366444
rect 70584 366392 70636 366444
rect 53472 366324 53524 366376
rect 171968 366324 172020 366376
rect 152464 365780 152516 365832
rect 276020 365780 276072 365832
rect 70584 365712 70636 365764
rect 291292 365712 291344 365764
rect 54852 365032 54904 365084
rect 96620 365032 96672 365084
rect 53748 364964 53800 365016
rect 202880 364964 202932 365016
rect 301044 364964 301096 365016
rect 96620 364420 96672 364472
rect 296904 364420 296956 364472
rect 158076 364352 158128 364404
rect 160744 364352 160796 364404
rect 179236 364352 179288 364404
rect 582380 364352 582432 364404
rect 160744 363740 160796 363792
rect 245844 363740 245896 363792
rect 162216 363672 162268 363724
rect 242808 363672 242860 363724
rect 347780 363672 347832 363724
rect 48044 363604 48096 363656
rect 62120 363604 62172 363656
rect 144184 363604 144236 363656
rect 178684 363604 178736 363656
rect 179328 363604 179380 363656
rect 580908 363604 580960 363656
rect 62120 362924 62172 362976
rect 62764 362924 62816 362976
rect 237472 362924 237524 362976
rect 240048 362924 240100 362976
rect 310520 362924 310572 362976
rect 287704 362312 287756 362364
rect 295432 362312 295484 362364
rect 55128 362176 55180 362228
rect 100760 362176 100812 362228
rect 171784 361632 171836 361684
rect 295524 361632 295576 361684
rect 100760 361564 100812 361616
rect 298284 361564 298336 361616
rect 122748 360816 122800 360868
rect 242900 360816 242952 360868
rect 250536 360408 250588 360460
rect 309784 360408 309836 360460
rect 187424 360340 187476 360392
rect 312544 360340 312596 360392
rect 31576 360272 31628 360324
rect 302332 360272 302384 360324
rect 171876 360204 171928 360256
rect 580264 360204 580316 360256
rect 163504 359456 163556 359508
rect 193864 359456 193916 359508
rect 166908 358980 166960 359032
rect 197728 358980 197780 359032
rect 172060 358912 172112 358964
rect 220084 358912 220136 358964
rect 220268 358912 220320 358964
rect 129096 358844 129148 358896
rect 202144 358844 202196 358896
rect 225420 358844 225472 358896
rect 302240 358844 302292 358896
rect 181628 358776 181680 358828
rect 337384 358776 337436 358828
rect 3332 358708 3384 358760
rect 17224 358708 17276 358760
rect 260104 358708 260156 358760
rect 266636 358708 266688 358760
rect 290464 357756 290516 357808
rect 308404 357756 308456 357808
rect 155868 357688 155920 357740
rect 182916 357688 182968 357740
rect 282092 357688 282144 357740
rect 313372 357688 313424 357740
rect 160008 357620 160060 357672
rect 184940 357620 184992 357672
rect 260748 357620 260800 357672
rect 305184 357620 305236 357672
rect 178776 357552 178828 357604
rect 211804 357552 211856 357604
rect 223488 357552 223540 357604
rect 298100 357552 298152 357604
rect 178684 357484 178736 357536
rect 218336 357484 218388 357536
rect 227352 357484 227404 357536
rect 342260 357484 342312 357536
rect 174636 357416 174688 357468
rect 262220 357416 262272 357468
rect 279424 357416 279476 357468
rect 449164 357416 449216 357468
rect 109040 357144 109092 357196
rect 109684 357144 109736 357196
rect 55128 356668 55180 356720
rect 80060 356668 80112 356720
rect 193220 356736 193272 356788
rect 109684 356668 109736 356720
rect 254216 356668 254268 356720
rect 289084 356668 289136 356720
rect 306472 356668 306524 356720
rect 171968 356260 172020 356312
rect 199660 356260 199712 356312
rect 174544 356192 174596 356244
rect 247132 356192 247184 356244
rect 247960 356192 248012 356244
rect 258908 356192 258960 356244
rect 294236 356192 294288 356244
rect 117964 356124 118016 356176
rect 214564 356124 214616 356176
rect 231124 356124 231176 356176
rect 345664 356124 345716 356176
rect 46756 356056 46808 356108
rect 305276 356056 305328 356108
rect 58992 355308 59044 355360
rect 131120 355308 131172 355360
rect 194600 355240 194652 355292
rect 195474 355240 195526 355292
rect 131120 355036 131172 355088
rect 283380 355036 283432 355088
rect 165436 354968 165488 355020
rect 209964 354968 210016 355020
rect 256976 354968 257028 355020
rect 297364 354968 297416 355020
rect 179880 354900 179932 354952
rect 287152 354900 287204 354952
rect 300124 354900 300176 354952
rect 170404 354832 170456 354884
rect 279056 354832 279108 354884
rect 285956 354832 286008 354884
rect 300952 354832 301004 354884
rect 68928 354764 68980 354816
rect 194600 354764 194652 354816
rect 269028 354764 269080 354816
rect 331496 354764 331548 354816
rect 275652 354696 275704 354748
rect 305092 354696 305144 354748
rect 292304 354492 292356 354544
rect 293316 354492 293368 354544
rect 175188 354356 175240 354408
rect 176660 354356 176712 354408
rect 170864 352656 170916 352708
rect 179788 352656 179840 352708
rect 90456 352588 90508 352640
rect 178776 352588 178828 352640
rect 49424 352520 49476 352572
rect 175188 352520 175240 352572
rect 175188 351908 175240 351960
rect 177580 351908 177632 351960
rect 52092 351160 52144 351212
rect 172060 351160 172112 351212
rect 50988 349800 51040 349852
rect 152556 349800 152608 349852
rect 63408 348372 63460 348424
rect 133972 348372 134024 348424
rect 134616 348372 134668 348424
rect 134616 347760 134668 347812
rect 176660 347760 176712 347812
rect 14464 347012 14516 347064
rect 35164 347012 35216 347064
rect 158628 345720 158680 345772
rect 176660 345720 176712 345772
rect 3332 345652 3384 345704
rect 14464 345652 14516 345704
rect 83464 345652 83516 345704
rect 171784 345652 171836 345704
rect 295616 345652 295668 345704
rect 468484 345652 468536 345704
rect 296076 343612 296128 343664
rect 296720 343612 296772 343664
rect 126888 341504 126940 341556
rect 179236 341504 179288 341556
rect 179512 341504 179564 341556
rect 132500 340892 132552 340944
rect 132868 340892 132920 340944
rect 160744 340892 160796 340944
rect 75920 340144 75972 340196
rect 132868 340144 132920 340196
rect 295616 339464 295668 339516
rect 309876 339464 309928 339516
rect 295616 339124 295668 339176
rect 298284 339124 298336 339176
rect 95056 338920 95108 338972
rect 102784 338920 102836 338972
rect 163596 333956 163648 334008
rect 176660 333956 176712 334008
rect 134524 333208 134576 333260
rect 176476 333208 176528 333260
rect 157248 329808 157300 329860
rect 176660 329808 176712 329860
rect 88340 329060 88392 329112
rect 162216 329060 162268 329112
rect 295524 327700 295576 327752
rect 347044 327700 347096 327752
rect 139492 327088 139544 327140
rect 176660 327088 176712 327140
rect 325056 324300 325108 324352
rect 580172 324300 580224 324352
rect 82728 323552 82780 323604
rect 106280 323552 106332 323604
rect 66076 322192 66128 322244
rect 164884 322192 164936 322244
rect 106280 321512 106332 321564
rect 163596 321512 163648 321564
rect 295432 320152 295484 320204
rect 336004 320152 336056 320204
rect 130476 319404 130528 319456
rect 162124 319404 162176 319456
rect 3424 319064 3476 319116
rect 8944 319064 8996 319116
rect 295432 318792 295484 318844
rect 350540 318792 350592 318844
rect 100668 318112 100720 318164
rect 133880 318112 133932 318164
rect 79324 318044 79376 318096
rect 158076 318044 158128 318096
rect 295432 317364 295484 317416
rect 302332 317364 302384 317416
rect 31576 316684 31628 316736
rect 70492 316684 70544 316736
rect 302332 316684 302384 316736
rect 467104 316684 467156 316736
rect 175096 316412 175148 316464
rect 177580 316412 177632 316464
rect 73160 315936 73212 315988
rect 169024 316004 169076 316056
rect 162768 315256 162820 315308
rect 176660 315256 176712 315308
rect 71872 314644 71924 314696
rect 73160 314644 73212 314696
rect 103612 314032 103664 314084
rect 134524 314032 134576 314084
rect 49608 313964 49660 314016
rect 126428 313964 126480 314016
rect 14464 313896 14516 313948
rect 118700 313896 118752 313948
rect 293868 313284 293920 313336
rect 356704 313284 356756 313336
rect 167736 313216 167788 313268
rect 170956 313216 171008 313268
rect 176660 313216 176712 313268
rect 300124 313216 300176 313268
rect 580172 313216 580224 313268
rect 8944 311788 8996 311840
rect 41420 311788 41472 311840
rect 50804 311176 50856 311228
rect 124312 311176 124364 311228
rect 41420 311108 41472 311160
rect 42616 311108 42668 311160
rect 116676 311108 116728 311160
rect 295340 310428 295392 310480
rect 305276 310428 305328 310480
rect 305460 310428 305512 310480
rect 116768 309816 116820 309868
rect 176660 309816 176712 309868
rect 41236 309748 41288 309800
rect 121552 309748 121604 309800
rect 305460 309748 305512 309800
rect 355324 309748 355376 309800
rect 43996 308456 44048 308508
rect 132500 308456 132552 308508
rect 33048 308388 33100 308440
rect 127808 308388 127860 308440
rect 295524 308388 295576 308440
rect 302332 308388 302384 308440
rect 98000 308116 98052 308168
rect 98736 308116 98788 308168
rect 98736 307776 98788 307828
rect 153936 307776 153988 307828
rect 81440 307368 81492 307420
rect 82084 307368 82136 307420
rect 75184 306416 75236 306468
rect 133144 306416 133196 306468
rect 81440 306348 81492 306400
rect 142896 306348 142948 306400
rect 68284 305668 68336 305720
rect 97264 305668 97316 305720
rect 46756 305600 46808 305652
rect 80060 305600 80112 305652
rect 121368 305600 121420 305652
rect 177856 305600 177908 305652
rect 86408 305056 86460 305108
rect 131856 305056 131908 305108
rect 3240 304988 3292 305040
rect 120080 304988 120132 305040
rect 121368 304988 121420 305040
rect 68836 304240 68888 304292
rect 174636 304240 174688 304292
rect 157156 303696 157208 303748
rect 176660 303696 176712 303748
rect 114008 303628 114060 303680
rect 171784 303628 171836 303680
rect 73804 303560 73856 303612
rect 88984 303560 89036 303612
rect 111800 302948 111852 303000
rect 132592 302948 132644 303000
rect 46848 302880 46900 302932
rect 69480 302880 69532 302932
rect 92388 302880 92440 302932
rect 115296 302880 115348 302932
rect 92848 302336 92900 302388
rect 162124 302336 162176 302388
rect 59084 302268 59136 302320
rect 145564 302268 145616 302320
rect 145748 302268 145800 302320
rect 69112 302200 69164 302252
rect 69480 302200 69532 302252
rect 167644 302200 167696 302252
rect 110880 301520 110932 301572
rect 111708 301520 111760 301572
rect 143632 301520 143684 301572
rect 91100 301452 91152 301504
rect 167736 301452 167788 301504
rect 97264 300840 97316 300892
rect 151084 300840 151136 300892
rect 295340 300840 295392 300892
rect 305276 300840 305328 300892
rect 142160 300772 142212 300824
rect 143448 300772 143500 300824
rect 94136 300568 94188 300620
rect 95148 300568 95200 300620
rect 108304 299820 108356 299872
rect 111800 299820 111852 299872
rect 84200 299752 84252 299804
rect 142988 299752 143040 299804
rect 95148 299684 95200 299736
rect 155316 299684 155368 299736
rect 79232 299616 79284 299668
rect 159456 299616 159508 299668
rect 77392 299548 77444 299600
rect 160836 299548 160888 299600
rect 32404 299480 32456 299532
rect 117964 299480 118016 299532
rect 143448 299480 143500 299532
rect 174636 299480 174688 299532
rect 167000 299412 167052 299464
rect 168288 299412 168340 299464
rect 176660 299412 176712 299464
rect 297364 299412 297416 299464
rect 580172 299412 580224 299464
rect 60464 298800 60516 298852
rect 120172 298800 120224 298852
rect 53564 298732 53616 298784
rect 167000 298732 167052 298784
rect 91744 298324 91796 298376
rect 133236 298324 133288 298376
rect 106740 298256 106792 298308
rect 148416 298256 148468 298308
rect 83556 298188 83608 298240
rect 145564 298188 145616 298240
rect 66168 298120 66220 298172
rect 140136 298120 140188 298172
rect 115940 298052 115992 298104
rect 116584 298052 116636 298104
rect 8208 297440 8260 297492
rect 72608 297440 72660 297492
rect 95056 297440 95108 297492
rect 176660 297440 176712 297492
rect 43904 297372 43956 297424
rect 129280 297372 129332 297424
rect 102232 296828 102284 296880
rect 148508 296828 148560 296880
rect 90640 296760 90692 296812
rect 138664 296760 138716 296812
rect 86132 296692 86184 296744
rect 151176 296692 151228 296744
rect 115112 295672 115164 295724
rect 116768 295672 116820 295724
rect 100944 295604 100996 295656
rect 127624 295604 127676 295656
rect 88064 295536 88116 295588
rect 126336 295536 126388 295588
rect 87420 295468 87472 295520
rect 131764 295468 131816 295520
rect 43444 295400 43496 295452
rect 100760 295400 100812 295452
rect 101588 295400 101640 295452
rect 110604 295400 110656 295452
rect 149980 295400 150032 295452
rect 82268 295332 82320 295384
rect 149796 295332 149848 295384
rect 295524 295332 295576 295384
rect 300124 295332 300176 295384
rect 50896 295264 50948 295316
rect 71780 295264 71832 295316
rect 174636 295264 174688 295316
rect 176660 295264 176712 295316
rect 64144 294584 64196 294636
rect 64696 294584 64748 294636
rect 70676 294584 70728 294636
rect 73252 294584 73304 294636
rect 75184 294584 75236 294636
rect 95792 294584 95844 294636
rect 173716 294584 173768 294636
rect 74540 294516 74592 294568
rect 91744 294516 91796 294568
rect 89812 294176 89864 294228
rect 95884 294176 95936 294228
rect 96436 294176 96488 294228
rect 105452 294176 105504 294228
rect 115940 294176 115992 294228
rect 123668 294176 123720 294228
rect 60004 294108 60056 294160
rect 92480 294108 92532 294160
rect 93860 294108 93912 294160
rect 124956 294108 125008 294160
rect 4804 293972 4856 294024
rect 79048 294040 79100 294092
rect 79324 294040 79376 294092
rect 80980 294040 81032 294092
rect 117964 294040 118016 294092
rect 77116 293972 77168 294024
rect 83464 293972 83516 294024
rect 85488 293972 85540 294024
rect 90456 293972 90508 294024
rect 91928 293972 91980 294024
rect 140044 293972 140096 294024
rect 295340 293972 295392 294024
rect 307024 293972 307076 294024
rect 103612 293904 103664 293956
rect 104532 293904 104584 293956
rect 109040 293904 109092 293956
rect 109684 293904 109736 293956
rect 46848 293292 46900 293344
rect 69020 293292 69072 293344
rect 2688 293224 2740 293276
rect 89812 293224 89864 293276
rect 98368 293224 98420 293276
rect 98644 293224 98696 293276
rect 68836 293088 68888 293140
rect 68836 292884 68888 292936
rect 116676 292884 116728 292936
rect 126520 292884 126572 292936
rect 92480 292816 92532 292868
rect 123760 292816 123812 292868
rect 99656 292748 99708 292800
rect 157984 292748 158036 292800
rect 75184 292680 75236 292732
rect 136088 292680 136140 292732
rect 58624 292612 58676 292664
rect 96712 292612 96764 292664
rect 98368 292612 98420 292664
rect 174636 292612 174688 292664
rect 69204 292544 69256 292596
rect 71964 292544 72016 292596
rect 84844 292544 84896 292596
rect 176016 292544 176068 292596
rect 67456 291864 67508 291916
rect 73712 291864 73764 291916
rect 83280 291864 83332 291916
rect 2872 291388 2924 291440
rect 8944 291388 8996 291440
rect 103152 291864 103204 291916
rect 112812 291864 112864 291916
rect 117320 291864 117372 291916
rect 120816 291864 120868 291916
rect 127716 291796 127768 291848
rect 143448 291796 143500 291848
rect 163596 291796 163648 291848
rect 137376 291320 137428 291372
rect 134616 291252 134668 291304
rect 129188 291184 129240 291236
rect 295616 291184 295668 291236
rect 301228 291184 301280 291236
rect 167000 291116 167052 291168
rect 168196 291116 168248 291168
rect 176660 291116 176712 291168
rect 295524 291116 295576 291168
rect 301044 291116 301096 291168
rect 17224 290436 17276 290488
rect 35808 290436 35860 290488
rect 52460 290436 52512 290488
rect 121460 289960 121512 290012
rect 144276 289960 144328 290012
rect 52460 289892 52512 289944
rect 53656 289892 53708 289944
rect 67732 289892 67784 289944
rect 121644 289892 121696 289944
rect 149888 289892 149940 289944
rect 48044 289824 48096 289876
rect 67640 289824 67692 289876
rect 121460 289756 121512 289808
rect 126428 289756 126480 289808
rect 172152 289824 172204 289876
rect 35808 289076 35860 289128
rect 67732 289076 67784 289128
rect 49608 288396 49660 288448
rect 67640 288396 67692 288448
rect 67456 288328 67508 288380
rect 67732 288328 67784 288380
rect 121460 288328 121512 288380
rect 170404 288328 170456 288380
rect 172428 288328 172480 288380
rect 176660 288328 176712 288380
rect 126428 287648 126480 287700
rect 139400 287648 139452 287700
rect 50896 287036 50948 287088
rect 67640 287036 67692 287088
rect 121644 287036 121696 287088
rect 155224 287036 155276 287088
rect 131212 285744 131264 285796
rect 132408 285744 132460 285796
rect 169392 285744 169444 285796
rect 54852 285676 54904 285728
rect 67824 285676 67876 285728
rect 124404 285676 124456 285728
rect 167920 285676 167972 285728
rect 295432 285676 295484 285728
rect 308588 285676 308640 285728
rect 121552 285608 121604 285660
rect 138020 285608 138072 285660
rect 121460 285540 121512 285592
rect 131212 285540 131264 285592
rect 122196 284928 122248 284980
rect 122840 284928 122892 284980
rect 130568 284928 130620 284980
rect 156604 284928 156656 284980
rect 43996 284316 44048 284368
rect 67640 284316 67692 284368
rect 53840 284248 53892 284300
rect 67732 284248 67784 284300
rect 160836 284248 160888 284300
rect 176660 284248 176712 284300
rect 66168 284180 66220 284232
rect 67640 284180 67692 284232
rect 295432 283568 295484 283620
rect 306564 283568 306616 283620
rect 325056 283568 325108 283620
rect 121460 282888 121512 282940
rect 173256 282888 173308 282940
rect 123760 282820 123812 282872
rect 166816 282820 166868 282872
rect 176660 282820 176712 282872
rect 121552 281596 121604 281648
rect 152556 281596 152608 281648
rect 32956 281528 33008 281580
rect 35716 281528 35768 281580
rect 121460 281528 121512 281580
rect 170404 281528 170456 281580
rect 295432 281528 295484 281580
rect 359464 281528 359516 281580
rect 67640 281460 67692 281512
rect 123668 280780 123720 280832
rect 160100 280780 160152 280832
rect 55036 280168 55088 280220
rect 67640 280168 67692 280220
rect 121460 280168 121512 280220
rect 136180 280168 136232 280220
rect 53748 280100 53800 280152
rect 67732 280100 67784 280152
rect 169116 280100 169168 280152
rect 176752 280100 176804 280152
rect 59084 280032 59136 280084
rect 67640 280032 67692 280084
rect 22744 279420 22796 279472
rect 59084 279420 59136 279472
rect 122748 279420 122800 279472
rect 173164 279420 173216 279472
rect 295432 278808 295484 278860
rect 297364 278808 297416 278860
rect 41236 278740 41288 278792
rect 57244 278740 57296 278792
rect 121460 278740 121512 278792
rect 141424 278740 141476 278792
rect 67640 278672 67692 278724
rect 121552 278672 121604 278724
rect 129740 278672 129792 278724
rect 160100 278060 160152 278112
rect 161388 278060 161440 278112
rect 176660 278060 176712 278112
rect 129740 277992 129792 278044
rect 131028 277992 131080 278044
rect 169208 277992 169260 278044
rect 52184 277380 52236 277432
rect 67640 277380 67692 277432
rect 121460 277312 121512 277364
rect 127808 277312 127860 277364
rect 145656 277380 145708 277432
rect 62028 276088 62080 276140
rect 64604 276088 64656 276140
rect 67640 276088 67692 276140
rect 50804 276020 50856 276072
rect 67732 276020 67784 276072
rect 295432 276020 295484 276072
rect 302424 276020 302476 276072
rect 306380 276020 306432 276072
rect 126520 275952 126572 276004
rect 176660 275952 176712 276004
rect 65524 275476 65576 275528
rect 68192 275476 68244 275528
rect 121460 274728 121512 274780
rect 148600 274728 148652 274780
rect 49516 274660 49568 274712
rect 67640 274660 67692 274712
rect 121552 274660 121604 274712
rect 164976 274660 165028 274712
rect 295432 274660 295484 274712
rect 301136 274660 301188 274712
rect 39948 274592 40000 274644
rect 68008 274592 68060 274644
rect 121460 274592 121512 274644
rect 179880 274592 179932 274644
rect 65984 273232 66036 273284
rect 67824 273232 67876 273284
rect 121460 273232 121512 273284
rect 158076 273232 158128 273284
rect 295432 272688 295484 272740
rect 298284 272688 298336 272740
rect 121460 272552 121512 272604
rect 124220 272552 124272 272604
rect 147128 272552 147180 272604
rect 128360 272484 128412 272536
rect 129280 272484 129332 272536
rect 176660 272484 176712 272536
rect 66168 271940 66220 271992
rect 67824 271940 67876 271992
rect 57796 271872 57848 271924
rect 67640 271872 67692 271924
rect 61844 270580 61896 270632
rect 67640 270580 67692 270632
rect 56324 270512 56376 270564
rect 67732 270512 67784 270564
rect 121460 270512 121512 270564
rect 138756 270512 138808 270564
rect 54944 269764 54996 269816
rect 67640 269764 67692 269816
rect 120908 269764 120960 269816
rect 128360 269764 128412 269816
rect 121460 269152 121512 269204
rect 154028 269152 154080 269204
rect 62028 269084 62080 269136
rect 67732 269084 67784 269136
rect 121552 269084 121604 269136
rect 160836 269084 160888 269136
rect 295432 269084 295484 269136
rect 349344 269084 349396 269136
rect 121460 269016 121512 269068
rect 135996 269016 136048 269068
rect 121460 268336 121512 268388
rect 126244 268336 126296 268388
rect 64788 267792 64840 267844
rect 67732 267792 67784 267844
rect 46756 267724 46808 267776
rect 67640 267724 67692 267776
rect 121552 267656 121604 267708
rect 148324 267656 148376 267708
rect 3424 266976 3476 267028
rect 13084 266976 13136 267028
rect 121460 266364 121512 266416
rect 166356 266364 166408 266416
rect 49424 266296 49476 266348
rect 67640 266296 67692 266348
rect 53472 264936 53524 264988
rect 68100 264936 68152 264988
rect 295432 264936 295484 264988
rect 325056 264936 325108 264988
rect 121460 264188 121512 264240
rect 159364 264188 159416 264240
rect 18604 263576 18656 263628
rect 59084 263576 59136 263628
rect 67640 263576 67692 263628
rect 121552 263576 121604 263628
rect 146944 263576 146996 263628
rect 121460 263508 121512 263560
rect 129832 263508 129884 263560
rect 4068 262828 4120 262880
rect 62120 262828 62172 262880
rect 121460 262828 121512 262880
rect 124312 262828 124364 262880
rect 140228 262828 140280 262880
rect 63316 262284 63368 262336
rect 67732 262284 67784 262336
rect 53748 262216 53800 262268
rect 67640 262216 67692 262268
rect 120724 262216 120776 262268
rect 121000 262216 121052 262268
rect 167736 262216 167788 262268
rect 62212 262148 62264 262200
rect 63040 262148 63092 262200
rect 67732 262148 67784 262200
rect 121460 262148 121512 262200
rect 171968 262148 172020 262200
rect 140136 262080 140188 262132
rect 176660 262080 176712 262132
rect 61752 261536 61804 261588
rect 61936 261536 61988 261588
rect 67640 261536 67692 261588
rect 50712 261468 50764 261520
rect 62212 261468 62264 261520
rect 52276 260856 52328 260908
rect 295432 260856 295484 260908
rect 309692 260856 309744 260908
rect 55864 260788 55916 260840
rect 67732 260788 67784 260840
rect 121460 260788 121512 260840
rect 161480 260788 161532 260840
rect 62120 260720 62172 260772
rect 67640 260720 67692 260772
rect 122104 260108 122156 260160
rect 141608 260108 141660 260160
rect 121460 259428 121512 259480
rect 160928 259428 160980 259480
rect 347044 259360 347096 259412
rect 580172 259360 580224 259412
rect 122288 258680 122340 258732
rect 171968 258680 172020 258732
rect 57704 258136 57756 258188
rect 67640 258136 67692 258188
rect 56416 258068 56468 258120
rect 67732 258068 67784 258120
rect 121460 258068 121512 258120
rect 162308 258068 162360 258120
rect 52092 258000 52144 258052
rect 67640 258000 67692 258052
rect 14464 257320 14516 257372
rect 52092 257320 52144 257372
rect 170956 257320 171008 257372
rect 178684 257320 178736 257372
rect 121552 256844 121604 256896
rect 148324 256844 148376 256896
rect 121460 256776 121512 256828
rect 156604 256776 156656 256828
rect 123576 256708 123628 256760
rect 176660 256708 176712 256760
rect 59268 255960 59320 256012
rect 67916 255960 67968 256012
rect 122472 255960 122524 256012
rect 130384 255960 130436 256012
rect 121552 255348 121604 255400
rect 135168 255348 135220 255400
rect 140780 255348 140832 255400
rect 60556 255280 60608 255332
rect 67640 255280 67692 255332
rect 121460 255280 121512 255332
rect 162400 255280 162452 255332
rect 41328 255212 41380 255264
rect 62120 255212 62172 255264
rect 62120 254532 62172 254584
rect 63132 254532 63184 254584
rect 67640 254532 67692 254584
rect 121460 253988 121512 254040
rect 151268 253988 151320 254040
rect 3424 253920 3476 253972
rect 26884 253920 26936 253972
rect 61936 253920 61988 253972
rect 67732 253920 67784 253972
rect 120724 253920 120776 253972
rect 172336 253920 172388 253972
rect 176660 253920 176712 253972
rect 295524 253920 295576 253972
rect 311164 253920 311216 253972
rect 62120 253852 62172 253904
rect 62764 253852 62816 253904
rect 67640 253852 67692 253904
rect 121460 253852 121512 253904
rect 166264 253852 166316 253904
rect 21364 253172 21416 253224
rect 62120 253172 62172 253224
rect 121552 252560 121604 252612
rect 138848 252560 138900 252612
rect 166724 252560 166776 252612
rect 176660 252560 176712 252612
rect 62120 251812 62172 251864
rect 63408 251812 63460 251864
rect 67640 251812 67692 251864
rect 295524 251812 295576 251864
rect 298376 251812 298428 251864
rect 305000 251812 305052 251864
rect 45192 251200 45244 251252
rect 62120 251200 62172 251252
rect 121460 251200 121512 251252
rect 176108 251200 176160 251252
rect 120632 251132 120684 251184
rect 133972 251132 134024 251184
rect 58716 249840 58768 249892
rect 67640 249840 67692 249892
rect 121552 249772 121604 249824
rect 134524 249772 134576 249824
rect 166816 249772 166868 249824
rect 176660 249772 176712 249824
rect 295524 249772 295576 249824
rect 325148 249772 325200 249824
rect 45468 249704 45520 249756
rect 67640 249704 67692 249756
rect 121460 249704 121512 249756
rect 130476 249704 130528 249756
rect 48228 249636 48280 249688
rect 58716 249636 58768 249688
rect 63132 248412 63184 248464
rect 67640 248412 67692 248464
rect 121460 248344 121512 248396
rect 174544 248344 174596 248396
rect 64696 247120 64748 247172
rect 67640 247120 67692 247172
rect 63224 247052 63276 247104
rect 67732 247052 67784 247104
rect 121552 247052 121604 247104
rect 144368 247052 144420 247104
rect 50988 246984 51040 247036
rect 67640 246984 67692 247036
rect 128360 246984 128412 247036
rect 132500 246984 132552 247036
rect 176660 246984 176712 247036
rect 66076 246916 66128 246968
rect 68192 246916 68244 246968
rect 139308 245760 139360 245812
rect 140136 245760 140188 245812
rect 121552 245692 121604 245744
rect 147036 245692 147088 245744
rect 121460 245624 121512 245676
rect 152648 245624 152700 245676
rect 295524 245624 295576 245676
rect 512644 245624 512696 245676
rect 121552 245556 121604 245608
rect 164240 245556 164292 245608
rect 121460 245012 121512 245064
rect 140136 245012 140188 245064
rect 134616 244944 134668 244996
rect 164884 244944 164936 244996
rect 120816 244876 120868 244928
rect 172060 244876 172112 244928
rect 66076 244264 66128 244316
rect 68192 244264 68244 244316
rect 8944 244196 8996 244248
rect 39672 244196 39724 244248
rect 67640 244196 67692 244248
rect 121460 244196 121512 244248
rect 153844 244196 153896 244248
rect 296904 242904 296956 242956
rect 347044 242904 347096 242956
rect 34428 242836 34480 242888
rect 69664 242836 69716 242888
rect 121552 242836 121604 242888
rect 143540 242836 143592 242888
rect 64604 242768 64656 242820
rect 66996 242768 67048 242820
rect 121460 242768 121512 242820
rect 127716 242768 127768 242820
rect 119988 242224 120040 242276
rect 155960 242224 156012 242276
rect 119896 242156 119948 242208
rect 179420 242156 179472 242208
rect 63408 241544 63460 241596
rect 67640 241544 67692 241596
rect 60464 241476 60516 241528
rect 67732 241476 67784 241528
rect 53564 241408 53616 241460
rect 67640 241408 67692 241460
rect 155316 241408 155368 241460
rect 298284 241408 298336 241460
rect 42708 240728 42760 240780
rect 63592 240728 63644 240780
rect 135168 240728 135220 240780
rect 190000 240592 190052 240644
rect 292028 240592 292080 240644
rect 293316 240592 293368 240644
rect 63592 240116 63644 240168
rect 64604 240116 64656 240168
rect 67640 240116 67692 240168
rect 121460 240116 121512 240168
rect 153844 240116 153896 240168
rect 163596 240048 163648 240100
rect 580172 240048 580224 240100
rect 121552 239980 121604 240032
rect 309140 239980 309192 240032
rect 310428 239980 310480 240032
rect 66260 239912 66312 239964
rect 70676 239912 70728 239964
rect 118976 239912 119028 239964
rect 119896 239912 119948 239964
rect 156604 239912 156656 239964
rect 306564 239912 306616 239964
rect 117044 239844 117096 239896
rect 120724 239844 120776 239896
rect 179420 239844 179472 239896
rect 301228 239844 301280 239896
rect 160744 239368 160796 239420
rect 168012 239368 168064 239420
rect 310428 239368 310480 239420
rect 331312 239368 331364 239420
rect 96436 239232 96488 239284
rect 97724 239232 97776 239284
rect 82912 239096 82964 239148
rect 292672 239096 292724 239148
rect 25504 239028 25556 239080
rect 81440 239028 81492 239080
rect 82268 239028 82320 239080
rect 63500 238960 63552 239012
rect 70032 238960 70084 239012
rect 107384 238960 107436 239012
rect 139492 238960 139544 239012
rect 48136 238892 48188 238944
rect 78680 238892 78732 238944
rect 79692 238892 79744 238944
rect 99380 238892 99432 238944
rect 99656 238892 99708 238944
rect 135904 238892 135956 238944
rect 59084 238824 59136 238876
rect 253020 238824 253072 238876
rect 298192 238824 298244 238876
rect 42524 238688 42576 238740
rect 82912 238688 82964 238740
rect 119804 238688 119856 238740
rect 124864 238688 124916 238740
rect 127532 238688 127584 238740
rect 250536 238688 250588 238740
rect 265532 238688 265584 238740
rect 299572 238688 299624 238740
rect 55128 238620 55180 238672
rect 89352 238620 89404 238672
rect 91928 238620 91980 238672
rect 149704 238620 149756 238672
rect 162308 238620 162360 238672
rect 276020 238620 276072 238672
rect 310612 238620 310664 238672
rect 59176 238552 59228 238604
rect 91284 238552 91336 238604
rect 105452 238552 105504 238604
rect 173808 238552 173860 238604
rect 176016 238552 176068 238604
rect 254400 238552 254452 238604
rect 288164 238552 288216 238604
rect 313280 238552 313332 238604
rect 99012 238484 99064 238536
rect 120908 238484 120960 238536
rect 169300 238484 169352 238536
rect 204904 238484 204956 238536
rect 240784 238484 240836 238536
rect 296076 238484 296128 238536
rect 117688 238416 117740 238468
rect 127532 238416 127584 238468
rect 174636 238416 174688 238468
rect 195980 238416 196032 238468
rect 88064 238348 88116 238400
rect 91744 238348 91796 238400
rect 108948 238348 109000 238400
rect 123484 238348 123536 238400
rect 96528 238280 96580 238332
rect 119896 238280 119948 238332
rect 60648 238144 60700 238196
rect 73068 238144 73120 238196
rect 73896 238144 73948 238196
rect 71320 238076 71372 238128
rect 86224 238076 86276 238128
rect 93216 238076 93268 238128
rect 98828 238076 98880 238128
rect 195980 238076 196032 238128
rect 210608 238076 210660 238128
rect 57888 238008 57940 238060
rect 92480 238008 92532 238060
rect 122288 238008 122340 238060
rect 327172 238008 327224 238060
rect 108028 237940 108080 237992
rect 108948 237940 109000 237992
rect 92480 237464 92532 237516
rect 93768 237464 93820 237516
rect 95148 237464 95200 237516
rect 70032 237396 70084 237448
rect 71044 237396 71096 237448
rect 75552 237396 75604 237448
rect 77116 237396 77168 237448
rect 2964 237328 3016 237380
rect 103520 237396 103572 237448
rect 104532 237396 104584 237448
rect 104624 237396 104676 237448
rect 106096 237396 106148 237448
rect 173808 237396 173860 237448
rect 175924 237396 175976 237448
rect 209320 237396 209372 237448
rect 210424 237396 210476 237448
rect 213184 237396 213236 237448
rect 216036 237396 216088 237448
rect 265624 237396 265676 237448
rect 267280 237396 267332 237448
rect 283564 237396 283616 237448
rect 284300 237396 284352 237448
rect 291936 237396 291988 237448
rect 292580 237396 292632 237448
rect 122472 237328 122524 237380
rect 322940 237328 322992 237380
rect 46664 237260 46716 237312
rect 106740 237260 106792 237312
rect 123576 237260 123628 237312
rect 145656 237260 145708 237312
rect 296904 237260 296956 237312
rect 45376 237192 45428 237244
rect 81624 237192 81676 237244
rect 95792 237192 95844 237244
rect 152464 237192 152516 237244
rect 162400 237192 162452 237244
rect 302424 237192 302476 237244
rect 41144 237124 41196 237176
rect 73252 237124 73304 237176
rect 98828 237124 98880 237176
rect 99288 237124 99340 237176
rect 126428 237124 126480 237176
rect 159364 237124 159416 237176
rect 269212 237124 269264 237176
rect 290464 237124 290516 237176
rect 300860 237124 300912 237176
rect 158168 237056 158220 237108
rect 191932 237056 191984 237108
rect 233884 237056 233936 237108
rect 299480 237056 299532 237108
rect 141516 236648 141568 236700
rect 239496 236648 239548 236700
rect 278780 236648 278832 236700
rect 294236 236648 294288 236700
rect 73252 235968 73304 236020
rect 73804 235968 73856 236020
rect 322940 235968 322992 236020
rect 323584 235968 323636 236020
rect 46756 235900 46808 235952
rect 302332 235900 302384 235952
rect 26884 235832 26936 235884
rect 112536 235832 112588 235884
rect 131120 235832 131172 235884
rect 176108 235832 176160 235884
rect 274088 235832 274140 235884
rect 306472 235832 306524 235884
rect 52368 235764 52420 235816
rect 80336 235764 80388 235816
rect 88248 235764 88300 235816
rect 126980 235764 127032 235816
rect 46848 235696 46900 235748
rect 71964 235696 72016 235748
rect 87420 235356 87472 235408
rect 88248 235356 88300 235408
rect 102232 235288 102284 235340
rect 129648 235356 129700 235408
rect 130568 235356 130620 235408
rect 166724 235356 166776 235408
rect 192484 235356 192536 235408
rect 151268 235288 151320 235340
rect 244924 235288 244976 235340
rect 60556 235220 60608 235272
rect 247684 235220 247736 235272
rect 250536 235220 250588 235272
rect 353944 235220 353996 235272
rect 46204 234608 46256 234660
rect 46756 234608 46808 234660
rect 71964 234608 72016 234660
rect 72424 234608 72476 234660
rect 80336 234608 80388 234660
rect 80704 234608 80756 234660
rect 56324 234540 56376 234592
rect 349252 234540 349304 234592
rect 63408 234472 63460 234524
rect 265532 234472 265584 234524
rect 13084 234404 13136 234456
rect 86868 234404 86920 234456
rect 110604 234404 110656 234456
rect 111064 234404 111116 234456
rect 129096 234404 129148 234456
rect 166356 234404 166408 234456
rect 317420 234472 317472 234524
rect 318064 234472 318116 234524
rect 83464 234336 83516 234388
rect 144184 234336 144236 234388
rect 160928 233996 160980 234048
rect 214564 233996 214616 234048
rect 171968 233928 172020 233980
rect 264336 233928 264388 233980
rect 84200 233860 84252 233912
rect 84844 233860 84896 233912
rect 89720 233860 89772 233912
rect 90640 233860 90692 233912
rect 93952 233860 94004 233912
rect 94504 233860 94556 233912
rect 100760 233860 100812 233912
rect 101588 233860 101640 233912
rect 103704 233860 103756 233912
rect 104808 233860 104860 233912
rect 114560 233860 114612 233912
rect 115756 233860 115808 233912
rect 169208 233860 169260 233912
rect 324596 233860 324648 233912
rect 114468 233248 114520 233300
rect 117964 233248 118016 233300
rect 61844 233180 61896 233232
rect 288164 233180 288216 233232
rect 347044 233180 347096 233232
rect 580172 233180 580224 233232
rect 113824 233112 113876 233164
rect 296812 233112 296864 233164
rect 45284 233044 45336 233096
rect 75184 233044 75236 233096
rect 75552 233044 75604 233096
rect 76472 233044 76524 233096
rect 137284 233044 137336 233096
rect 148600 233044 148652 233096
rect 295524 233044 295576 233096
rect 44088 232976 44140 233028
rect 77760 232976 77812 233028
rect 77944 232976 77996 233028
rect 86868 232976 86920 233028
rect 195980 232976 196032 233028
rect 27528 232908 27580 232960
rect 113180 232908 113232 232960
rect 114468 232908 114520 232960
rect 167920 232908 167972 232960
rect 271144 232908 271196 232960
rect 311164 232568 311216 232620
rect 335452 232568 335504 232620
rect 282184 232500 282236 232552
rect 313372 232500 313424 232552
rect 128360 231820 128412 231872
rect 129004 231820 129056 231872
rect 346584 231820 346636 231872
rect 61936 231752 61988 231804
rect 298376 231752 298428 231804
rect 81624 231684 81676 231736
rect 278872 231684 278924 231736
rect 37096 231616 37148 231668
rect 104256 231616 104308 231668
rect 104624 231616 104676 231668
rect 169760 231616 169812 231668
rect 171048 231616 171100 231668
rect 305276 231616 305328 231668
rect 115112 231548 115164 231600
rect 179788 231548 179840 231600
rect 236000 231548 236052 231600
rect 88708 231480 88760 231532
rect 128360 231480 128412 231532
rect 154488 231140 154540 231192
rect 169760 231140 169812 231192
rect 173256 231140 173308 231192
rect 222844 231140 222896 231192
rect 68744 231072 68796 231124
rect 325792 231072 325844 231124
rect 39764 230392 39816 230444
rect 104164 230392 104216 230444
rect 104532 230392 104584 230444
rect 154488 230392 154540 230444
rect 172060 230392 172112 230444
rect 332600 230392 332652 230444
rect 98368 230324 98420 230376
rect 233884 230324 233936 230376
rect 118332 230256 118384 230308
rect 240784 230256 240836 230308
rect 63224 229780 63276 229832
rect 161480 229780 161532 229832
rect 161388 229712 161440 229764
rect 574744 229712 574796 229764
rect 74724 229032 74776 229084
rect 294144 229032 294196 229084
rect 38568 228964 38620 229016
rect 122932 228964 122984 229016
rect 155224 228964 155276 229016
rect 328552 228964 328604 229016
rect 69112 228896 69164 228948
rect 241520 228896 241572 228948
rect 159456 228352 159508 228404
rect 255320 228352 255372 228404
rect 122932 227740 122984 227792
rect 124864 227740 124916 227792
rect 53656 227672 53708 227724
rect 287704 227672 287756 227724
rect 108672 227604 108724 227656
rect 153108 227604 153160 227656
rect 163504 227604 163556 227656
rect 218060 227604 218112 227656
rect 145564 227196 145616 227248
rect 232504 227196 232556 227248
rect 100944 227128 100996 227180
rect 198188 227128 198240 227180
rect 60464 227060 60516 227112
rect 158168 227060 158220 227112
rect 231860 227060 231912 227112
rect 268384 227060 268436 227112
rect 153108 226992 153160 227044
rect 329932 226992 329984 227044
rect 63316 226244 63368 226296
rect 290464 226244 290516 226296
rect 177672 225632 177724 225684
rect 189724 225632 189776 225684
rect 148324 225564 148376 225616
rect 240784 225564 240836 225616
rect 325056 225564 325108 225616
rect 332600 225564 332652 225616
rect 81440 224884 81492 224936
rect 277400 224884 277452 224936
rect 3424 224204 3476 224256
rect 120172 224204 120224 224256
rect 136180 224204 136232 224256
rect 239404 224204 239456 224256
rect 68836 223524 68888 223576
rect 324320 223524 324372 223576
rect 140228 222912 140280 222964
rect 287796 222912 287848 222964
rect 79048 222844 79100 222896
rect 273260 222844 273312 222896
rect 325148 222844 325200 222896
rect 333980 222844 334032 222896
rect 170404 221484 170456 221536
rect 203524 221484 203576 221536
rect 64604 221416 64656 221468
rect 343640 221416 343692 221468
rect 58716 220192 58768 220244
rect 122104 220192 122156 220244
rect 141608 220192 141660 220244
rect 283656 220192 283708 220244
rect 89996 220124 90048 220176
rect 252836 220124 252888 220176
rect 65984 220056 66036 220108
rect 251180 220056 251232 220108
rect 256700 220056 256752 220108
rect 278044 220056 278096 220108
rect 239496 219376 239548 219428
rect 327080 219376 327132 219428
rect 335360 219376 335412 219428
rect 355324 219376 355376 219428
rect 580172 219376 580224 219428
rect 52276 218900 52328 218952
rect 163504 218900 163556 218952
rect 164976 218900 165028 218952
rect 269120 218900 269172 218952
rect 99472 218832 99524 218884
rect 220084 218832 220136 218884
rect 142896 218764 142948 218816
rect 307116 218764 307168 218816
rect 50712 218696 50764 218748
rect 311164 218696 311216 218748
rect 55036 217404 55088 217456
rect 196716 217404 196768 217456
rect 67548 217336 67600 217388
rect 251272 217336 251324 217388
rect 71044 217268 71096 217320
rect 315396 217268 315448 217320
rect 122196 216588 122248 216640
rect 304264 216656 304316 216708
rect 346676 216656 346728 216708
rect 93952 216520 94004 216572
rect 146300 216520 146352 216572
rect 142988 216112 143040 216164
rect 235264 216112 235316 216164
rect 50896 216044 50948 216096
rect 162308 216044 162360 216096
rect 146300 215976 146352 216028
rect 327080 215976 327132 216028
rect 74632 215908 74684 215960
rect 280160 215908 280212 215960
rect 258080 215364 258132 215416
rect 264244 215364 264296 215416
rect 3332 215228 3384 215280
rect 18604 215228 18656 215280
rect 103704 215228 103756 215280
rect 164148 215228 164200 215280
rect 154028 214820 154080 214872
rect 270592 214820 270644 214872
rect 50804 214752 50856 214804
rect 211804 214752 211856 214804
rect 164148 214684 164200 214736
rect 328460 214684 328512 214736
rect 57796 214616 57848 214668
rect 250444 214616 250496 214668
rect 108948 214548 109000 214600
rect 328644 214548 328696 214600
rect 84292 213868 84344 213920
rect 133880 213868 133932 213920
rect 135168 213868 135220 213920
rect 147036 213324 147088 213376
rect 259460 213324 259512 213376
rect 111800 213256 111852 213308
rect 273352 213256 273404 213308
rect 25504 213188 25556 213240
rect 83464 213188 83516 213240
rect 135168 213188 135220 213240
rect 322940 213188 322992 213240
rect 137376 211964 137428 212016
rect 224224 211964 224276 212016
rect 62028 211896 62080 211948
rect 272064 211896 272116 211948
rect 78680 211828 78732 211880
rect 328552 211828 328604 211880
rect 35716 211760 35768 211812
rect 313924 211760 313976 211812
rect 289820 211148 289872 211200
rect 296720 211148 296772 211200
rect 89720 210536 89772 210588
rect 253940 210536 253992 210588
rect 129648 210468 129700 210520
rect 335360 210468 335412 210520
rect 53472 210400 53524 210452
rect 289084 210400 289136 210452
rect 43996 209720 44048 209772
rect 327264 209720 327316 209772
rect 84200 209652 84252 209704
rect 136640 209652 136692 209704
rect 126336 209176 126388 209228
rect 233884 209176 233936 209228
rect 136640 209108 136692 209160
rect 321652 209108 321704 209160
rect 86224 209040 86276 209092
rect 277400 209040 277452 209092
rect 327264 209040 327316 209092
rect 354680 209040 354732 209092
rect 114560 208292 114612 208344
rect 169760 208292 169812 208344
rect 80060 208224 80112 208276
rect 122840 208224 122892 208276
rect 124128 208224 124180 208276
rect 169760 207884 169812 207936
rect 170864 207884 170916 207936
rect 186964 207884 187016 207936
rect 158076 207816 158128 207868
rect 233976 207816 234028 207868
rect 245660 207816 245712 207868
rect 308496 207816 308548 207868
rect 115940 207748 115992 207800
rect 246304 207748 246356 207800
rect 124128 207680 124180 207732
rect 330116 207680 330168 207732
rect 54944 207612 54996 207664
rect 318156 207612 318208 207664
rect 574744 206932 574796 206984
rect 579896 206932 579948 206984
rect 248420 206592 248472 206644
rect 287704 206592 287756 206644
rect 149980 206524 150032 206576
rect 270684 206524 270736 206576
rect 168012 206456 168064 206508
rect 345020 206456 345072 206508
rect 66168 206388 66220 206440
rect 251364 206388 251416 206440
rect 274640 206388 274692 206440
rect 293224 206388 293276 206440
rect 133144 206320 133196 206372
rect 350632 206320 350684 206372
rect 104256 206252 104308 206304
rect 339592 206252 339644 206304
rect 96436 205572 96488 205624
rect 146208 205572 146260 205624
rect 146208 205028 146260 205080
rect 346492 205028 346544 205080
rect 48044 204960 48096 205012
rect 278964 204960 279016 205012
rect 74540 204892 74592 204944
rect 343732 204892 343784 204944
rect 146944 203804 146996 203856
rect 264980 203804 265032 203856
rect 133236 203736 133288 203788
rect 267832 203736 267884 203788
rect 110420 203668 110472 203720
rect 249800 203668 249852 203720
rect 271880 203668 271932 203720
rect 294052 203668 294104 203720
rect 92480 203600 92532 203652
rect 242164 203600 242216 203652
rect 281540 203600 281592 203652
rect 342352 203600 342404 203652
rect 72424 203532 72476 203584
rect 325884 203532 325936 203584
rect 119988 202240 120040 202292
rect 329840 202240 329892 202292
rect 66076 202172 66128 202224
rect 278872 202172 278924 202224
rect 99380 202104 99432 202156
rect 327356 202104 327408 202156
rect 158168 200880 158220 200932
rect 256976 200880 257028 200932
rect 131856 200812 131908 200864
rect 318248 200812 318300 200864
rect 153936 200744 153988 200796
rect 351920 200744 351972 200796
rect 157984 199588 158036 199640
rect 246396 199588 246448 199640
rect 134524 199520 134576 199572
rect 242256 199520 242308 199572
rect 69296 199452 69348 199504
rect 248512 199452 248564 199504
rect 93768 199384 93820 199436
rect 347872 199384 347924 199436
rect 160836 198160 160888 198212
rect 266360 198160 266412 198212
rect 138664 198092 138716 198144
rect 276112 198092 276164 198144
rect 126244 198024 126296 198076
rect 311256 198024 311308 198076
rect 77944 197956 77996 198008
rect 330024 197956 330076 198008
rect 144368 196868 144420 196920
rect 262404 196868 262456 196920
rect 222844 196800 222896 196852
rect 354772 196800 354824 196852
rect 96620 196732 96672 196784
rect 249064 196732 249116 196784
rect 63132 196664 63184 196716
rect 271972 196664 272024 196716
rect 56416 196596 56468 196648
rect 276020 196596 276072 196648
rect 138848 195440 138900 195492
rect 239496 195440 239548 195492
rect 91744 195372 91796 195424
rect 246488 195372 246540 195424
rect 163504 195304 163556 195356
rect 334256 195304 334308 195356
rect 160744 195236 160796 195288
rect 582472 195236 582524 195288
rect 99288 194012 99340 194064
rect 162400 194012 162452 194064
rect 124956 193944 125008 193996
rect 231124 193944 231176 193996
rect 144276 193876 144328 193928
rect 266452 193876 266504 193928
rect 140136 193808 140188 193860
rect 340972 193808 341024 193860
rect 227720 192720 227772 192772
rect 346400 192720 346452 192772
rect 100760 192652 100812 192704
rect 254032 192652 254084 192704
rect 77300 192584 77352 192636
rect 252652 192584 252704 192636
rect 104164 192516 104216 192568
rect 321560 192516 321612 192568
rect 49608 192448 49660 192500
rect 269212 192448 269264 192500
rect 124864 191360 124916 191412
rect 185584 191360 185636 191412
rect 204168 191360 204220 191412
rect 220820 191360 220872 191412
rect 136088 191292 136140 191344
rect 242348 191292 242400 191344
rect 148508 191224 148560 191276
rect 255412 191224 255464 191276
rect 53748 191156 53800 191208
rect 259552 191156 259604 191208
rect 264336 191156 264388 191208
rect 342536 191156 342588 191208
rect 70400 191088 70452 191140
rect 315488 191088 315540 191140
rect 214564 190068 214616 190120
rect 274824 190068 274876 190120
rect 160008 190000 160060 190052
rect 196624 190000 196676 190052
rect 237380 190000 237432 190052
rect 340880 190000 340932 190052
rect 153844 189932 153896 189984
rect 258172 189932 258224 189984
rect 102140 189864 102192 189916
rect 249984 189864 250036 189916
rect 18604 189796 18656 189848
rect 109040 189796 109092 189848
rect 169392 189796 169444 189848
rect 341064 189796 341116 189848
rect 88248 189728 88300 189780
rect 327264 189728 327316 189780
rect 106188 189116 106240 189168
rect 169208 189116 169260 189168
rect 134524 189048 134576 189100
rect 214656 189048 214708 189100
rect 3424 188980 3476 189032
rect 60004 188980 60056 189032
rect 140044 188436 140096 188488
rect 263692 188436 263744 188488
rect 127624 188368 127676 188420
rect 269304 188368 269356 188420
rect 66996 188300 67048 188352
rect 319536 188300 319588 188352
rect 102048 187688 102100 187740
rect 184204 187688 184256 187740
rect 157156 187212 157208 187264
rect 198096 187212 198148 187264
rect 131764 187144 131816 187196
rect 267740 187144 267792 187196
rect 173164 187076 173216 187128
rect 324504 187076 324556 187128
rect 49516 187008 49568 187060
rect 256792 187008 256844 187060
rect 96528 186940 96580 186992
rect 321836 186940 321888 186992
rect 323676 186940 323728 186992
rect 332692 186940 332744 186992
rect 132408 186396 132460 186448
rect 167920 186396 167972 186448
rect 104808 186328 104860 186380
rect 173256 186328 173308 186380
rect 196716 185784 196768 185836
rect 259644 185784 259696 185836
rect 141424 185716 141476 185768
rect 255596 185716 255648 185768
rect 148416 185648 148468 185700
rect 318432 185648 318484 185700
rect 73804 185580 73856 185632
rect 321284 185580 321336 185632
rect 100668 184968 100720 185020
rect 170404 184968 170456 185020
rect 125508 184900 125560 184952
rect 214932 184900 214984 184952
rect 155868 184492 155920 184544
rect 192576 184492 192628 184544
rect 203524 184492 203576 184544
rect 259736 184492 259788 184544
rect 149796 184424 149848 184476
rect 274732 184424 274784 184476
rect 64696 184356 64748 184408
rect 254216 184356 254268 184408
rect 319444 184356 319496 184408
rect 332784 184356 332836 184408
rect 111156 184288 111208 184340
rect 339776 184288 339828 184340
rect 69664 184220 69716 184272
rect 338396 184220 338448 184272
rect 75184 184152 75236 184204
rect 347964 184152 348016 184204
rect 157248 182996 157300 183048
rect 191104 182996 191156 183048
rect 224224 182996 224276 183048
rect 260932 182996 260984 183048
rect 162216 182928 162268 182980
rect 338212 182928 338264 182980
rect 122104 182860 122156 182912
rect 345204 182860 345256 182912
rect 73068 182792 73120 182844
rect 336832 182792 336884 182844
rect 118424 182180 118476 182232
rect 167828 182180 167880 182232
rect 240784 181704 240836 181756
rect 262220 181704 262272 181756
rect 232504 181636 232556 181688
rect 258264 181636 258316 181688
rect 318064 181636 318116 181688
rect 338304 181636 338356 181688
rect 94044 181568 94096 181620
rect 249892 181568 249944 181620
rect 289084 181568 289136 181620
rect 334072 181568 334124 181620
rect 167736 181500 167788 181552
rect 345112 181500 345164 181552
rect 41236 181432 41288 181484
rect 313832 181432 313884 181484
rect 314568 181432 314620 181484
rect 336740 181432 336792 181484
rect 133604 180888 133656 180940
rect 164332 180888 164384 180940
rect 122012 180820 122064 180872
rect 211988 180820 212040 180872
rect 244924 180344 244976 180396
rect 255504 180344 255556 180396
rect 242164 180276 242216 180328
rect 256884 180276 256936 180328
rect 244280 180208 244332 180260
rect 270500 180208 270552 180260
rect 167644 180140 167696 180192
rect 196716 180140 196768 180192
rect 233976 180140 234028 180192
rect 260840 180140 260892 180192
rect 64788 180072 64840 180124
rect 251456 180072 251508 180124
rect 315304 180072 315356 180124
rect 341156 180072 341208 180124
rect 123024 179596 123076 179648
rect 166356 179596 166408 179648
rect 121000 179528 121052 179580
rect 167736 179528 167788 179580
rect 128176 179460 128228 179512
rect 214104 179460 214156 179512
rect 114284 179392 114336 179444
rect 209044 179392 209096 179444
rect 172152 179324 172204 179376
rect 346308 179324 346360 179376
rect 169024 179256 169076 179308
rect 342628 179256 342680 179308
rect 242348 178780 242400 178832
rect 258448 178780 258500 178832
rect 211804 178712 211856 178764
rect 258080 178712 258132 178764
rect 311256 178712 311308 178764
rect 332692 178712 332744 178764
rect 138756 178644 138808 178696
rect 252560 178644 252612 178696
rect 312544 178644 312596 178696
rect 338120 178644 338172 178696
rect 112444 178236 112496 178288
rect 211896 178236 211948 178288
rect 130752 178168 130804 178220
rect 165528 178168 165580 178220
rect 148232 178100 148284 178152
rect 214564 178100 214616 178152
rect 159916 178032 159968 178084
rect 167644 178032 167696 178084
rect 289084 178032 289136 178084
rect 316040 178032 316092 178084
rect 52552 177964 52604 178016
rect 120080 177964 120132 178016
rect 242256 177964 242308 178016
rect 249340 177964 249392 178016
rect 109960 177896 110012 177948
rect 134524 177896 134576 177948
rect 239496 177556 239548 177608
rect 256700 177556 256752 177608
rect 246488 177488 246540 177540
rect 267924 177488 267976 177540
rect 315488 177488 315540 177540
rect 331404 177488 331456 177540
rect 233884 177420 233936 177472
rect 258356 177420 258408 177472
rect 311164 177420 311216 177472
rect 331220 177420 331272 177472
rect 220084 177352 220136 177404
rect 262312 177352 262364 177404
rect 289728 177352 289780 177404
rect 310520 177352 310572 177404
rect 313924 177352 313976 177404
rect 335544 177352 335596 177404
rect 166816 177284 166868 177336
rect 198004 177284 198056 177336
rect 198188 177284 198240 177336
rect 263600 177284 263652 177336
rect 287796 177284 287848 177336
rect 334164 177284 334216 177336
rect 134432 177012 134484 177064
rect 165252 177012 165304 177064
rect 127072 176944 127124 176996
rect 173164 176944 173216 176996
rect 125784 176876 125836 176928
rect 188344 176876 188396 176928
rect 108120 176808 108172 176860
rect 170496 176808 170548 176860
rect 107016 176740 107068 176792
rect 169300 176740 169352 176792
rect 135720 176672 135772 176724
rect 213920 176604 213972 176656
rect 235264 176604 235316 176656
rect 248052 176604 248104 176656
rect 313832 176604 313884 176656
rect 321468 176604 321520 176656
rect 319536 176536 319588 176588
rect 321744 176536 321796 176588
rect 129464 176264 129516 176316
rect 166172 176264 166224 176316
rect 119436 176196 119488 176248
rect 166448 176196 166500 176248
rect 115756 176128 115808 176180
rect 166264 176128 166316 176180
rect 98368 176060 98420 176112
rect 169024 176060 169076 176112
rect 100760 175992 100812 176044
rect 171876 175992 171928 176044
rect 13084 175924 13136 175976
rect 111064 175924 111116 175976
rect 116952 175924 117004 175976
rect 169116 175924 169168 175976
rect 246304 175924 246356 175976
rect 252744 175924 252796 175976
rect 315396 175924 315448 175976
rect 332876 175924 332928 175976
rect 166540 175244 166592 175296
rect 343824 175244 343876 175296
rect 165252 175176 165304 175228
rect 213920 175176 213972 175228
rect 164332 175108 164384 175160
rect 214012 175108 214064 175160
rect 2780 164092 2832 164144
rect 4804 164092 4856 164144
rect 3424 150356 3476 150408
rect 17224 150356 17276 150408
rect 3240 137912 3292 137964
rect 14464 137912 14516 137964
rect 63408 125604 63460 125656
rect 66168 125604 66220 125656
rect 63316 121456 63368 121508
rect 66076 121456 66128 121508
rect 3424 111732 3476 111784
rect 13084 111732 13136 111784
rect 3424 97928 3476 97980
rect 25504 97928 25556 97980
rect 262864 174496 262916 174548
rect 274088 174496 274140 174548
rect 287980 174020 288032 174072
rect 307576 174020 307628 174072
rect 271144 173952 271196 174004
rect 307300 173952 307352 174004
rect 265900 173884 265952 173936
rect 307668 173884 307720 173936
rect 165528 173816 165580 173868
rect 214012 173816 214064 173868
rect 252468 173816 252520 173868
rect 258080 173816 258132 173868
rect 167920 173748 167972 173800
rect 213920 173748 213972 173800
rect 258080 173680 258132 173732
rect 258356 173680 258408 173732
rect 251732 172796 251784 172848
rect 255596 172796 255648 172848
rect 283656 172660 283708 172712
rect 307576 172660 307628 172712
rect 269764 172592 269816 172644
rect 307300 172592 307352 172644
rect 265716 172524 265768 172576
rect 307668 172524 307720 172576
rect 166172 172456 166224 172508
rect 213920 172456 213972 172508
rect 252468 172388 252520 172440
rect 260840 172388 260892 172440
rect 252376 172320 252428 172372
rect 262404 172320 262456 172372
rect 281080 171164 281132 171216
rect 306932 171164 306984 171216
rect 262956 171096 263008 171148
rect 307484 171096 307536 171148
rect 173164 171028 173216 171080
rect 213920 171028 213972 171080
rect 188344 170960 188396 171012
rect 214012 170960 214064 171012
rect 324320 170892 324372 170944
rect 325976 170892 326028 170944
rect 251548 170756 251600 170808
rect 254216 170756 254268 170808
rect 169300 170348 169352 170400
rect 214840 170348 214892 170400
rect 252284 170280 252336 170332
rect 256792 170280 256844 170332
rect 304264 169872 304316 169924
rect 307484 169872 307536 169924
rect 273904 169804 273956 169856
rect 307300 169804 307352 169856
rect 267188 169736 267240 169788
rect 307668 169736 307720 169788
rect 166356 169668 166408 169720
rect 213920 169668 213972 169720
rect 324320 169668 324372 169720
rect 331220 169668 331272 169720
rect 252192 169600 252244 169652
rect 258080 169600 258132 169652
rect 170496 168988 170548 169040
rect 215024 168988 215076 169040
rect 287888 168512 287940 168564
rect 307668 168512 307720 168564
rect 279424 168444 279476 168496
rect 307576 168444 307628 168496
rect 264336 168376 264388 168428
rect 307300 168376 307352 168428
rect 167736 168308 167788 168360
rect 213920 168308 213972 168360
rect 252468 168308 252520 168360
rect 263692 168308 263744 168360
rect 324320 168308 324372 168360
rect 338396 168308 338448 168360
rect 211988 168240 212040 168292
rect 214012 168240 214064 168292
rect 294604 167696 294656 167748
rect 307024 167696 307076 167748
rect 258908 167628 258960 167680
rect 307392 167628 307444 167680
rect 252284 167424 252336 167476
rect 256700 167424 256752 167476
rect 267096 167016 267148 167068
rect 306932 167016 306984 167068
rect 166448 166948 166500 167000
rect 213920 166948 213972 167000
rect 167828 166880 167880 166932
rect 214012 166880 214064 166932
rect 169116 166812 169168 166864
rect 213920 166812 213972 166864
rect 252284 166812 252336 166864
rect 258172 166812 258224 166864
rect 251916 166404 251968 166456
rect 259552 166404 259604 166456
rect 249708 166268 249760 166320
rect 305184 166268 305236 166320
rect 252284 166064 252336 166116
rect 256884 166064 256936 166116
rect 282368 165724 282420 165776
rect 306932 165724 306984 165776
rect 272524 165656 272576 165708
rect 307484 165656 307536 165708
rect 257528 165588 257580 165640
rect 307668 165588 307720 165640
rect 166264 165520 166316 165572
rect 213920 165520 213972 165572
rect 252468 165520 252520 165572
rect 270684 165520 270736 165572
rect 324412 165520 324464 165572
rect 335360 165520 335412 165572
rect 209044 165452 209096 165504
rect 214012 165452 214064 165504
rect 324320 165452 324372 165504
rect 332876 165452 332928 165504
rect 251548 164432 251600 164484
rect 252836 164432 252888 164484
rect 278136 164364 278188 164416
rect 307668 164364 307720 164416
rect 271236 164296 271288 164348
rect 307576 164296 307628 164348
rect 260196 164228 260248 164280
rect 307300 164228 307352 164280
rect 211896 164160 211948 164212
rect 213920 164160 213972 164212
rect 252468 164160 252520 164212
rect 267832 164160 267884 164212
rect 324320 164160 324372 164212
rect 339776 164160 339828 164212
rect 252100 164092 252152 164144
rect 264980 164092 265032 164144
rect 324412 164092 324464 164144
rect 334256 164092 334308 164144
rect 261116 163480 261168 163532
rect 291844 163480 291896 163532
rect 290648 162936 290700 162988
rect 307300 162936 307352 162988
rect 268476 162868 268528 162920
rect 307668 162868 307720 162920
rect 252468 162800 252520 162852
rect 270592 162800 270644 162852
rect 324320 162800 324372 162852
rect 353300 162800 353352 162852
rect 263048 162120 263100 162172
rect 307208 162120 307260 162172
rect 252468 161916 252520 161968
rect 259644 161916 259696 161968
rect 298744 161508 298796 161560
rect 307484 161508 307536 161560
rect 258816 161440 258868 161492
rect 307668 161440 307720 161492
rect 324320 161372 324372 161424
rect 341064 161372 341116 161424
rect 252468 161032 252520 161084
rect 258264 161032 258316 161084
rect 252468 160896 252520 160948
rect 259736 160896 259788 160948
rect 167920 160760 167972 160812
rect 192668 160760 192720 160812
rect 177764 160692 177816 160744
rect 215944 160692 215996 160744
rect 261484 160692 261536 160744
rect 307116 160692 307168 160744
rect 302976 160216 303028 160268
rect 307668 160216 307720 160268
rect 283748 160148 283800 160200
rect 306748 160148 306800 160200
rect 253572 160080 253624 160132
rect 255320 160080 255372 160132
rect 260104 160080 260156 160132
rect 307484 160080 307536 160132
rect 169208 160012 169260 160064
rect 213920 160012 213972 160064
rect 252468 160012 252520 160064
rect 269212 160012 269264 160064
rect 324320 160012 324372 160064
rect 331404 160012 331456 160064
rect 173256 159944 173308 159996
rect 214012 159944 214064 159996
rect 251916 159944 251968 159996
rect 266452 159944 266504 159996
rect 259000 159332 259052 159384
rect 307392 159332 307444 159384
rect 301504 158788 301556 158840
rect 307668 158788 307720 158840
rect 265808 158720 265860 158772
rect 307576 158720 307628 158772
rect 184204 158652 184256 158704
rect 213920 158652 213972 158704
rect 324412 158652 324464 158704
rect 343916 158652 343968 158704
rect 324320 158584 324372 158636
rect 332784 158584 332836 158636
rect 252560 157972 252612 158024
rect 260932 157972 260984 158024
rect 296076 157496 296128 157548
rect 307668 157496 307720 157548
rect 264428 157428 264480 157480
rect 306932 157428 306984 157480
rect 257436 157360 257488 157412
rect 307300 157360 307352 157412
rect 170404 157292 170456 157344
rect 214012 157292 214064 157344
rect 251548 157292 251600 157344
rect 274824 157292 274876 157344
rect 324320 157292 324372 157344
rect 336924 157292 336976 157344
rect 171876 157224 171928 157276
rect 213920 157224 213972 157276
rect 252468 157224 252520 157276
rect 269304 157224 269356 157276
rect 324412 157156 324464 157208
rect 327356 157156 327408 157208
rect 278412 156612 278464 156664
rect 307668 156612 307720 156664
rect 269856 156000 269908 156052
rect 307484 156000 307536 156052
rect 261576 155932 261628 155984
rect 306748 155932 306800 155984
rect 169024 155864 169076 155916
rect 213920 155864 213972 155916
rect 252376 155864 252428 155916
rect 276112 155864 276164 155916
rect 324320 155864 324372 155916
rect 356060 155864 356112 155916
rect 252468 155796 252520 155848
rect 263600 155796 263652 155848
rect 204904 155184 204956 155236
rect 216128 155184 216180 155236
rect 251732 155184 251784 155236
rect 269120 155184 269172 155236
rect 285220 154708 285272 154760
rect 307576 154708 307628 154760
rect 276756 154640 276808 154692
rect 307668 154640 307720 154692
rect 253480 154572 253532 154624
rect 307484 154572 307536 154624
rect 252008 154504 252060 154556
rect 277400 154504 277452 154556
rect 324320 154504 324372 154556
rect 346584 154504 346636 154556
rect 251548 154436 251600 154488
rect 272064 154436 272116 154488
rect 324412 154436 324464 154488
rect 330116 154436 330168 154488
rect 252468 154368 252520 154420
rect 267924 154368 267976 154420
rect 282460 153824 282512 153876
rect 307392 153824 307444 153876
rect 204996 153280 205048 153332
rect 214012 153280 214064 153332
rect 269948 153280 270000 153332
rect 307668 153280 307720 153332
rect 202144 153212 202196 153264
rect 213920 153212 213972 153264
rect 261668 153212 261720 153264
rect 307484 153212 307536 153264
rect 252284 153144 252336 153196
rect 278964 153144 279016 153196
rect 324320 153144 324372 153196
rect 341156 153144 341208 153196
rect 250812 152668 250864 152720
rect 258356 152668 258408 152720
rect 250536 152600 250588 152652
rect 261024 152600 261076 152652
rect 251824 152532 251876 152584
rect 272524 152532 272576 152584
rect 255964 152464 256016 152516
rect 307576 152464 307628 152516
rect 195244 151852 195296 151904
rect 213920 151852 213972 151904
rect 285128 151852 285180 151904
rect 307484 151852 307536 151904
rect 184204 151784 184256 151836
rect 214012 151784 214064 151836
rect 275560 151784 275612 151836
rect 307668 151784 307720 151836
rect 324412 151716 324464 151768
rect 336832 151716 336884 151768
rect 252376 151648 252428 151700
rect 262312 151648 262364 151700
rect 324320 151648 324372 151700
rect 328644 151648 328696 151700
rect 252468 151580 252520 151632
rect 273352 151580 273404 151632
rect 251272 151240 251324 151292
rect 253940 151240 253992 151292
rect 177856 151036 177908 151088
rect 211804 151036 211856 151088
rect 256332 151036 256384 151088
rect 306656 151036 306708 151088
rect 274180 150492 274232 150544
rect 307484 150492 307536 150544
rect 206376 150424 206428 150476
rect 213920 150424 213972 150476
rect 258724 150424 258776 150476
rect 307668 150424 307720 150476
rect 192668 150356 192720 150408
rect 214012 150356 214064 150408
rect 252468 150356 252520 150408
rect 274732 150356 274784 150408
rect 324320 150356 324372 150408
rect 346676 150356 346728 150408
rect 254676 149676 254728 149728
rect 306564 149676 306616 149728
rect 251732 149608 251784 149660
rect 255504 149608 255556 149660
rect 303160 149200 303212 149252
rect 307300 149200 307352 149252
rect 276664 149132 276716 149184
rect 306932 149132 306984 149184
rect 260380 149064 260432 149116
rect 307484 149064 307536 149116
rect 167644 148996 167696 149048
rect 213920 148996 213972 149048
rect 252468 148996 252520 149048
rect 280160 148996 280212 149048
rect 324320 148996 324372 149048
rect 338304 148996 338356 149048
rect 251548 148384 251600 148436
rect 255412 148384 255464 148436
rect 254768 148316 254820 148368
rect 307208 148316 307260 148368
rect 252376 147704 252428 147756
rect 256976 147704 257028 147756
rect 272616 147704 272668 147756
rect 307484 147704 307536 147756
rect 185676 147636 185728 147688
rect 213920 147636 213972 147688
rect 257344 147636 257396 147688
rect 307668 147636 307720 147688
rect 252468 147568 252520 147620
rect 267740 147568 267792 147620
rect 324320 147568 324372 147620
rect 347780 147568 347832 147620
rect 251272 147228 251324 147280
rect 254032 147228 254084 147280
rect 177304 146888 177356 146940
rect 214104 146888 214156 146940
rect 284944 146412 284996 146464
rect 307668 146412 307720 146464
rect 256240 146344 256292 146396
rect 306748 146344 306800 146396
rect 203524 146276 203576 146328
rect 213920 146276 213972 146328
rect 256148 146276 256200 146328
rect 307576 146276 307628 146328
rect 252468 146208 252520 146260
rect 276020 146208 276072 146260
rect 252100 146140 252152 146192
rect 273260 146140 273312 146192
rect 261760 145528 261812 145580
rect 307024 145528 307076 145580
rect 211896 144984 211948 145036
rect 214472 144984 214524 145036
rect 299020 144984 299072 145036
rect 307484 144984 307536 145036
rect 170404 144916 170456 144968
rect 213920 144916 213972 144968
rect 254584 144916 254636 144968
rect 307668 144916 307720 144968
rect 252468 144848 252520 144900
rect 266360 144848 266412 144900
rect 324320 144848 324372 144900
rect 345204 144848 345256 144900
rect 252100 144780 252152 144832
rect 262220 144780 262272 144832
rect 299112 144168 299164 144220
rect 307300 144168 307352 144220
rect 251548 143624 251600 143676
rect 259460 143624 259512 143676
rect 279608 143624 279660 143676
rect 307484 143624 307536 143676
rect 167644 143556 167696 143608
rect 213920 143556 213972 143608
rect 253388 143556 253440 143608
rect 306932 143556 306984 143608
rect 324320 143488 324372 143540
rect 335544 143488 335596 143540
rect 251916 142808 251968 142860
rect 269856 142808 269908 142860
rect 301688 142264 301740 142316
rect 307392 142264 307444 142316
rect 271328 142196 271380 142248
rect 306748 142196 306800 142248
rect 209044 142128 209096 142180
rect 213920 142128 213972 142180
rect 253296 142128 253348 142180
rect 307668 142128 307720 142180
rect 252468 141924 252520 141976
rect 256792 141924 256844 141976
rect 262864 141380 262916 141432
rect 306564 141380 306616 141432
rect 304356 140904 304408 140956
rect 307668 140904 307720 140956
rect 289360 140836 289412 140888
rect 307576 140836 307628 140888
rect 182824 140768 182876 140820
rect 213920 140768 213972 140820
rect 275468 140768 275520 140820
rect 307484 140768 307536 140820
rect 251180 140428 251232 140480
rect 253572 140428 253624 140480
rect 184480 140020 184532 140072
rect 214656 140020 214708 140072
rect 193864 139476 193916 139528
rect 214012 139476 214064 139528
rect 181444 139408 181496 139460
rect 213920 139408 213972 139460
rect 280896 139408 280948 139460
rect 307668 139408 307720 139460
rect 252468 139340 252520 139392
rect 278872 139340 278924 139392
rect 324320 139340 324372 139392
rect 338212 139340 338264 139392
rect 468484 139340 468536 139392
rect 580172 139340 580224 139392
rect 251732 138728 251784 138780
rect 271144 138728 271196 138780
rect 250720 138660 250772 138712
rect 300952 138660 301004 138712
rect 297548 138116 297600 138168
rect 307668 138116 307720 138168
rect 207664 138048 207716 138100
rect 214012 138048 214064 138100
rect 290556 138048 290608 138100
rect 307576 138048 307628 138100
rect 192668 137980 192720 138032
rect 213920 137980 213972 138032
rect 272524 137980 272576 138032
rect 307484 137980 307536 138032
rect 252468 137912 252520 137964
rect 271972 137912 272024 137964
rect 324320 137912 324372 137964
rect 345112 137912 345164 137964
rect 324504 137844 324556 137896
rect 328552 137844 328604 137896
rect 251272 137708 251324 137760
rect 254124 137708 254176 137760
rect 323584 137300 323636 137352
rect 324412 137300 324464 137352
rect 187056 137232 187108 137284
rect 214472 137232 214524 137284
rect 267004 136756 267056 136808
rect 307484 136756 307536 136808
rect 250628 136688 250680 136740
rect 307576 136688 307628 136740
rect 169116 136620 169168 136672
rect 214104 136620 214156 136672
rect 250444 136620 250496 136672
rect 307668 136620 307720 136672
rect 252468 136552 252520 136604
rect 294604 136552 294656 136604
rect 252100 136484 252152 136536
rect 265900 136484 265952 136536
rect 252192 135940 252244 135992
rect 278136 135940 278188 135992
rect 264888 135872 264940 135924
rect 302240 135872 302292 135924
rect 302884 135396 302936 135448
rect 307484 135396 307536 135448
rect 172060 135328 172112 135380
rect 214012 135328 214064 135380
rect 294696 135328 294748 135380
rect 307668 135328 307720 135380
rect 169024 135260 169076 135312
rect 213920 135260 213972 135312
rect 278320 135260 278372 135312
rect 306932 135260 306984 135312
rect 252468 135192 252520 135244
rect 283656 135192 283708 135244
rect 324320 135192 324372 135244
rect 350632 135192 350684 135244
rect 252284 135124 252336 135176
rect 269764 135124 269816 135176
rect 324504 135124 324556 135176
rect 342444 135124 342496 135176
rect 269948 134512 270000 134564
rect 307300 134512 307352 134564
rect 279516 134036 279568 134088
rect 307484 134036 307536 134088
rect 295984 133968 296036 134020
rect 307668 133968 307720 134020
rect 166264 133900 166316 133952
rect 213920 133900 213972 133952
rect 251272 133832 251324 133884
rect 281080 133832 281132 133884
rect 324320 133832 324372 133884
rect 331312 133832 331364 133884
rect 252468 133764 252520 133816
rect 265716 133764 265768 133816
rect 252376 133696 252428 133748
rect 262956 133696 263008 133748
rect 280804 133220 280856 133272
rect 298100 133220 298152 133272
rect 263140 133152 263192 133204
rect 307116 133152 307168 133204
rect 301596 132608 301648 132660
rect 307668 132608 307720 132660
rect 282276 132540 282328 132592
rect 306932 132540 306984 132592
rect 173164 132472 173216 132524
rect 213920 132472 213972 132524
rect 280988 132472 281040 132524
rect 306564 132472 306616 132524
rect 251732 132404 251784 132456
rect 304264 132404 304316 132456
rect 324320 132404 324372 132456
rect 354772 132404 354824 132456
rect 252284 132336 252336 132388
rect 258908 132336 258960 132388
rect 252008 131724 252060 131776
rect 285128 131724 285180 131776
rect 285036 131180 285088 131232
rect 307668 131180 307720 131232
rect 283840 131112 283892 131164
rect 306932 131112 306984 131164
rect 252284 131044 252336 131096
rect 279424 131044 279476 131096
rect 324320 131044 324372 131096
rect 343824 131044 343876 131096
rect 252376 130976 252428 131028
rect 273904 130976 273956 131028
rect 252468 130908 252520 130960
rect 267188 130908 267240 130960
rect 256700 130364 256752 130416
rect 305092 130364 305144 130416
rect 174544 129820 174596 129872
rect 213920 129820 213972 129872
rect 278228 129820 278280 129872
rect 307300 129820 307352 129872
rect 171876 129752 171928 129804
rect 214012 129752 214064 129804
rect 273996 129752 274048 129804
rect 307668 129752 307720 129804
rect 252468 129684 252520 129736
rect 287888 129684 287940 129736
rect 324412 129684 324464 129736
rect 329840 129684 329892 129736
rect 252376 129616 252428 129668
rect 264336 129616 264388 129668
rect 324320 129616 324372 129668
rect 330024 129616 330076 129668
rect 252284 129548 252336 129600
rect 261484 129548 261536 129600
rect 287796 128460 287848 128512
rect 307668 128460 307720 128512
rect 286324 128392 286376 128444
rect 307300 128392 307352 128444
rect 188344 128324 188396 128376
rect 213920 128324 213972 128376
rect 269856 128324 269908 128376
rect 306748 128324 306800 128376
rect 251824 128256 251876 128308
rect 282368 128256 282420 128308
rect 324412 128256 324464 128308
rect 347964 128256 348016 128308
rect 252468 128188 252520 128240
rect 267096 128188 267148 128240
rect 324320 128188 324372 128240
rect 329932 128188 329984 128240
rect 252376 128120 252428 128172
rect 263048 128120 263100 128172
rect 171784 127576 171836 127628
rect 210608 127576 210660 127628
rect 294788 127576 294840 127628
rect 307208 127576 307260 127628
rect 189816 127032 189868 127084
rect 213920 127032 213972 127084
rect 279424 127032 279476 127084
rect 307576 127032 307628 127084
rect 171968 126964 172020 127016
rect 214012 126964 214064 127016
rect 271144 126964 271196 127016
rect 307668 126964 307720 127016
rect 252192 126896 252244 126948
rect 271236 126896 271288 126948
rect 324320 126896 324372 126948
rect 342536 126896 342588 126948
rect 449164 126896 449216 126948
rect 580172 126896 580224 126948
rect 252468 126692 252520 126744
rect 257528 126692 257580 126744
rect 276020 126284 276072 126336
rect 292028 126284 292080 126336
rect 251548 126216 251600 126268
rect 305644 126216 305696 126268
rect 211988 125672 212040 125724
rect 214748 125672 214800 125724
rect 289176 125672 289228 125724
rect 306564 125672 306616 125724
rect 166356 125604 166408 125656
rect 213920 125604 213972 125656
rect 260288 125604 260340 125656
rect 306932 125604 306984 125656
rect 252468 125060 252520 125112
rect 259000 125060 259052 125112
rect 252192 124856 252244 124908
rect 301504 124856 301556 124908
rect 252468 124584 252520 124636
rect 260196 124584 260248 124636
rect 264336 124380 264388 124432
rect 306932 124380 306984 124432
rect 184388 124244 184440 124296
rect 214012 124244 214064 124296
rect 265716 124244 265768 124296
rect 307668 124244 307720 124296
rect 167736 124176 167788 124228
rect 213920 124176 213972 124228
rect 301780 124176 301832 124228
rect 307484 124176 307536 124228
rect 252468 124108 252520 124160
rect 290648 124108 290700 124160
rect 324320 124108 324372 124160
rect 334164 124108 334216 124160
rect 251272 124040 251324 124092
rect 268476 124040 268528 124092
rect 251824 123428 251876 123480
rect 284944 123428 284996 123480
rect 290464 122952 290516 123004
rect 307576 122952 307628 123004
rect 176016 122884 176068 122936
rect 214012 122884 214064 122936
rect 287888 122884 287940 122936
rect 307668 122884 307720 122936
rect 170496 122816 170548 122868
rect 213920 122816 213972 122868
rect 285128 122816 285180 122868
rect 307484 122816 307536 122868
rect 252468 122748 252520 122800
rect 298744 122748 298796 122800
rect 324320 122748 324372 122800
rect 351920 122748 351972 122800
rect 252376 122680 252428 122732
rect 261760 122680 261812 122732
rect 324412 122680 324464 122732
rect 343732 122680 343784 122732
rect 251732 122612 251784 122664
rect 258816 122612 258868 122664
rect 173348 122068 173400 122120
rect 214748 122068 214800 122120
rect 300216 121592 300268 121644
rect 307484 121592 307536 121644
rect 210516 121524 210568 121576
rect 214012 121524 214064 121576
rect 283656 121524 283708 121576
rect 307668 121524 307720 121576
rect 188436 121456 188488 121508
rect 213920 121456 213972 121508
rect 261484 121456 261536 121508
rect 306932 121456 306984 121508
rect 252376 121388 252428 121440
rect 302976 121388 303028 121440
rect 324412 121388 324464 121440
rect 339684 121388 339736 121440
rect 252468 121320 252520 121372
rect 283748 121320 283800 121372
rect 251732 121252 251784 121304
rect 260104 121252 260156 121304
rect 324320 120980 324372 121032
rect 327080 120980 327132 121032
rect 171784 120708 171836 120760
rect 214932 120708 214984 120760
rect 304540 120232 304592 120284
rect 307484 120232 307536 120284
rect 298928 120164 298980 120216
rect 306748 120164 306800 120216
rect 196808 120096 196860 120148
rect 213920 120096 213972 120148
rect 273904 120096 273956 120148
rect 307668 120096 307720 120148
rect 252284 120028 252336 120080
rect 265808 120028 265860 120080
rect 324320 120028 324372 120080
rect 340972 120028 341024 120080
rect 251456 119960 251508 120012
rect 254768 119960 254820 120012
rect 252100 119824 252152 119876
rect 260380 119824 260432 119876
rect 260104 119348 260156 119400
rect 307024 119348 307076 119400
rect 182916 118804 182968 118856
rect 213920 118804 213972 118856
rect 301504 118804 301556 118856
rect 306564 118804 306616 118856
rect 177488 118736 177540 118788
rect 214012 118736 214064 118788
rect 293224 118736 293276 118788
rect 307668 118736 307720 118788
rect 166448 118668 166500 118720
rect 214104 118668 214156 118720
rect 269764 118668 269816 118720
rect 306932 118668 306984 118720
rect 251732 118600 251784 118652
rect 296076 118600 296128 118652
rect 324412 118600 324464 118652
rect 347872 118600 347924 118652
rect 252468 118532 252520 118584
rect 264428 118532 264480 118584
rect 324320 118532 324372 118584
rect 339592 118532 339644 118584
rect 264980 117920 265032 117972
rect 293132 117920 293184 117972
rect 252284 117852 252336 117904
rect 257436 117852 257488 117904
rect 302976 117444 303028 117496
rect 307576 117444 307628 117496
rect 185768 117376 185820 117428
rect 214012 117376 214064 117428
rect 297456 117376 297508 117428
rect 307668 117376 307720 117428
rect 167828 117308 167880 117360
rect 213920 117308 213972 117360
rect 292028 117308 292080 117360
rect 306564 117308 306616 117360
rect 251272 117240 251324 117292
rect 278412 117240 278464 117292
rect 252468 117172 252520 117224
rect 261576 117172 261628 117224
rect 282368 116084 282420 116136
rect 307668 116084 307720 116136
rect 169300 116016 169352 116068
rect 214012 116016 214064 116068
rect 278136 116016 278188 116068
rect 306748 116016 306800 116068
rect 169208 115948 169260 116000
rect 213920 115948 213972 116000
rect 262956 115948 263008 116000
rect 307576 115948 307628 116000
rect 251548 115880 251600 115932
rect 282460 115880 282512 115932
rect 324412 115880 324464 115932
rect 354680 115880 354732 115932
rect 324320 115812 324372 115864
rect 336740 115812 336792 115864
rect 251180 115608 251232 115660
rect 253480 115608 253532 115660
rect 304448 114656 304500 114708
rect 306748 114656 306800 114708
rect 203616 114588 203668 114640
rect 214012 114588 214064 114640
rect 297640 114588 297692 114640
rect 307576 114588 307628 114640
rect 173256 114520 173308 114572
rect 213920 114520 213972 114572
rect 268476 114520 268528 114572
rect 307668 114520 307720 114572
rect 252468 114452 252520 114504
rect 285220 114452 285272 114504
rect 324320 114452 324372 114504
rect 346492 114452 346544 114504
rect 252376 114384 252428 114436
rect 276756 114384 276808 114436
rect 324412 114384 324464 114436
rect 343640 114384 343692 114436
rect 252468 114316 252520 114368
rect 261668 114316 261720 114368
rect 170772 113772 170824 113824
rect 199384 113772 199436 113824
rect 177396 113228 177448 113280
rect 213920 113228 213972 113280
rect 294604 113228 294656 113280
rect 307668 113228 307720 113280
rect 170588 113160 170640 113212
rect 214012 113160 214064 113212
rect 284944 113160 284996 113212
rect 307576 113160 307628 113212
rect 324320 113092 324372 113144
rect 332692 113092 332744 113144
rect 467104 113092 467156 113144
rect 579804 113092 579856 113144
rect 251732 112956 251784 113008
rect 255964 112956 256016 113008
rect 252100 112616 252152 112668
rect 256332 112616 256384 112668
rect 252376 112412 252428 112464
rect 299020 112412 299072 112464
rect 300308 111936 300360 111988
rect 307668 111936 307720 111988
rect 207756 111868 207808 111920
rect 214012 111868 214064 111920
rect 298836 111868 298888 111920
rect 307484 111868 307536 111920
rect 189908 111800 189960 111852
rect 213920 111800 213972 111852
rect 256056 111800 256108 111852
rect 307576 111800 307628 111852
rect 167920 111732 167972 111784
rect 206376 111732 206428 111784
rect 252100 111732 252152 111784
rect 275560 111732 275612 111784
rect 324320 111732 324372 111784
rect 345020 111732 345072 111784
rect 324412 111664 324464 111716
rect 334072 111664 334124 111716
rect 251640 111392 251692 111444
rect 254676 111392 254728 111444
rect 251916 111052 251968 111104
rect 279608 111052 279660 111104
rect 304264 110576 304316 110628
rect 307668 110576 307720 110628
rect 200764 110508 200816 110560
rect 214012 110508 214064 110560
rect 283748 110508 283800 110560
rect 307484 110508 307536 110560
rect 184296 110440 184348 110492
rect 213920 110440 213972 110492
rect 275376 110440 275428 110492
rect 307576 110440 307628 110492
rect 168104 110372 168156 110424
rect 177304 110372 177356 110424
rect 252100 110372 252152 110424
rect 301688 110372 301740 110424
rect 324320 110372 324372 110424
rect 339500 110372 339552 110424
rect 251548 110304 251600 110356
rect 274180 110304 274232 110356
rect 252468 109488 252520 109540
rect 258724 109488 258776 109540
rect 304356 109148 304408 109200
rect 307484 109148 307536 109200
rect 178684 109080 178736 109132
rect 214012 109080 214064 109132
rect 299020 109080 299072 109132
rect 307576 109080 307628 109132
rect 168012 109012 168064 109064
rect 213920 109012 213972 109064
rect 271236 109012 271288 109064
rect 307668 109012 307720 109064
rect 167920 108944 167972 108996
rect 184480 108944 184532 108996
rect 252008 108944 252060 108996
rect 303160 108944 303212 108996
rect 252468 108876 252520 108928
rect 276664 108876 276716 108928
rect 267096 107856 267148 107908
rect 307668 107856 307720 107908
rect 205088 107720 205140 107772
rect 213920 107720 213972 107772
rect 300400 107720 300452 107772
rect 307576 107720 307628 107772
rect 188528 107652 188580 107704
rect 214012 107652 214064 107704
rect 303068 107652 303120 107704
rect 306932 107652 306984 107704
rect 251824 107584 251876 107636
rect 272616 107584 272668 107636
rect 252100 107516 252152 107568
rect 263140 107516 263192 107568
rect 252468 107448 252520 107500
rect 257344 107448 257396 107500
rect 301688 106428 301740 106480
rect 307484 106428 307536 106480
rect 192760 106360 192812 106412
rect 213920 106360 213972 106412
rect 276664 106360 276716 106412
rect 307576 106360 307628 106412
rect 174636 106292 174688 106344
rect 214012 106292 214064 106344
rect 261576 106292 261628 106344
rect 307668 106292 307720 106344
rect 252008 106224 252060 106276
rect 299112 106224 299164 106276
rect 252284 106088 252336 106140
rect 254584 106088 254636 106140
rect 252468 105748 252520 105800
rect 256240 105748 256292 105800
rect 255964 105544 256016 105596
rect 295340 105544 295392 105596
rect 212080 105000 212132 105052
rect 214104 105000 214156 105052
rect 296076 105000 296128 105052
rect 307484 105000 307536 105052
rect 206468 104932 206520 104984
rect 213920 104932 213972 104984
rect 298744 104932 298796 104984
rect 307668 104932 307720 104984
rect 194048 104864 194100 104916
rect 214012 104864 214064 104916
rect 252468 104796 252520 104848
rect 294788 104796 294840 104848
rect 324320 104796 324372 104848
rect 328460 104796 328512 104848
rect 252192 104660 252244 104712
rect 256148 104660 256200 104712
rect 251364 104116 251416 104168
rect 287980 104116 288032 104168
rect 303160 103640 303212 103692
rect 307576 103640 307628 103692
rect 206376 103572 206428 103624
rect 214012 103572 214064 103624
rect 294880 103572 294932 103624
rect 307668 103572 307720 103624
rect 177304 103504 177356 103556
rect 213920 103504 213972 103556
rect 293316 103504 293368 103556
rect 307484 103504 307536 103556
rect 252468 103436 252520 103488
rect 262864 103436 262916 103488
rect 324320 103300 324372 103352
rect 327264 103300 327316 103352
rect 170956 102756 171008 102808
rect 204904 102756 204956 102808
rect 251180 102756 251232 102808
rect 253388 102756 253440 102808
rect 251272 102688 251324 102740
rect 293960 102756 294012 102808
rect 296168 102280 296220 102332
rect 306748 102280 306800 102332
rect 294788 102212 294840 102264
rect 307668 102212 307720 102264
rect 209228 102144 209280 102196
rect 213920 102144 213972 102196
rect 261668 102144 261720 102196
rect 307484 102144 307536 102196
rect 252468 102076 252520 102128
rect 271328 102076 271380 102128
rect 324320 102076 324372 102128
rect 349252 102076 349304 102128
rect 251180 101940 251232 101992
rect 253296 101940 253348 101992
rect 170680 101396 170732 101448
rect 214656 101396 214708 101448
rect 252192 101396 252244 101448
rect 289084 101396 289136 101448
rect 292120 100784 292172 100836
rect 306564 100784 306616 100836
rect 173440 100716 173492 100768
rect 213920 100716 213972 100768
rect 250536 100716 250588 100768
rect 307668 100716 307720 100768
rect 252008 100648 252060 100700
rect 289360 100648 289412 100700
rect 512644 100648 512696 100700
rect 580172 100648 580224 100700
rect 252468 100580 252520 100632
rect 275468 100580 275520 100632
rect 251548 100512 251600 100564
rect 269948 100512 270000 100564
rect 209136 99424 209188 99476
rect 214012 99424 214064 99476
rect 289268 99424 289320 99476
rect 307576 99424 307628 99476
rect 164884 99356 164936 99408
rect 213920 99356 213972 99408
rect 274180 99356 274232 99408
rect 307668 99356 307720 99408
rect 252468 98812 252520 98864
rect 260104 98812 260156 98864
rect 293408 98132 293460 98184
rect 307668 98132 307720 98184
rect 187148 98064 187200 98116
rect 213920 98064 213972 98116
rect 260196 98064 260248 98116
rect 307484 98064 307536 98116
rect 166540 97996 166592 98048
rect 214012 97996 214064 98048
rect 256148 97996 256200 98048
rect 307576 97996 307628 98048
rect 251180 97928 251232 97980
rect 253204 97928 253256 97980
rect 289084 96772 289136 96824
rect 306748 96772 306800 96824
rect 262864 96704 262916 96756
rect 307668 96704 307720 96756
rect 193956 96636 194008 96688
rect 213920 96636 213972 96688
rect 253296 96636 253348 96688
rect 307484 96636 307536 96688
rect 258080 95888 258132 95940
rect 283564 95888 283616 95940
rect 318064 95752 318116 95804
rect 321468 95752 321520 95804
rect 185584 95140 185636 95192
rect 323124 95140 323176 95192
rect 186964 95072 187016 95124
rect 321652 95072 321704 95124
rect 199384 95004 199436 95056
rect 321744 95004 321796 95056
rect 131948 94120 132000 94172
rect 170404 94120 170456 94172
rect 151912 94052 151964 94104
rect 195244 94052 195296 94104
rect 151728 93984 151780 94036
rect 204996 93984 205048 94036
rect 109040 93916 109092 93968
rect 169300 93916 169352 93968
rect 113732 93848 113784 93900
rect 177488 93848 177540 93900
rect 241520 93848 241572 93900
rect 250720 93848 250772 93900
rect 175924 93780 175976 93832
rect 324504 93780 324556 93832
rect 63316 93712 63368 93764
rect 209228 93712 209280 93764
rect 210608 93712 210660 93764
rect 321560 93712 321612 93764
rect 64788 93644 64840 93696
rect 206468 93644 206520 93696
rect 121736 93304 121788 93356
rect 176016 93304 176068 93356
rect 124496 93236 124548 93288
rect 182824 93236 182876 93288
rect 107752 93168 107804 93220
rect 169208 93168 169260 93220
rect 102048 93100 102100 93152
rect 174544 93100 174596 93152
rect 119344 92420 119396 92472
rect 207664 92420 207716 92472
rect 120356 92352 120408 92404
rect 181444 92352 181496 92404
rect 115480 92284 115532 92336
rect 170680 92284 170732 92336
rect 133144 92216 133196 92268
rect 187056 92216 187108 92268
rect 151728 92148 151780 92200
rect 202144 92148 202196 92200
rect 125968 92080 126020 92132
rect 171784 92080 171836 92132
rect 228364 91876 228416 91928
rect 260288 91876 260340 91928
rect 192576 91808 192628 91860
rect 232504 91808 232556 91860
rect 179144 91740 179196 91792
rect 245660 91740 245712 91792
rect 94228 91264 94280 91316
rect 120724 91264 120776 91316
rect 101864 91196 101916 91248
rect 127624 91196 127676 91248
rect 85948 91128 86000 91180
rect 120816 91128 120868 91180
rect 74816 91060 74868 91112
rect 112444 91060 112496 91112
rect 67364 90992 67416 91044
rect 214932 90992 214984 91044
rect 66168 90924 66220 90976
rect 177304 90924 177356 90976
rect 196716 90924 196768 90976
rect 323032 90924 323084 90976
rect 124128 90856 124180 90908
rect 184388 90856 184440 90908
rect 115204 90788 115256 90840
rect 166448 90788 166500 90840
rect 122840 90720 122892 90772
rect 167736 90720 167788 90772
rect 151728 90652 151780 90704
rect 184204 90652 184256 90704
rect 309692 90380 309744 90432
rect 320180 90380 320232 90432
rect 308588 90312 308640 90364
rect 328460 90312 328512 90364
rect 89076 89632 89128 89684
rect 209136 89632 209188 89684
rect 123944 89564 123996 89616
rect 213184 89564 213236 89616
rect 112352 89496 112404 89548
rect 182916 89496 182968 89548
rect 104532 89428 104584 89480
rect 170588 89428 170640 89480
rect 106924 89360 106976 89412
rect 173164 89360 173216 89412
rect 126612 89292 126664 89344
rect 166356 89292 166408 89344
rect 91008 88272 91060 88324
rect 212080 88272 212132 88324
rect 106648 88204 106700 88256
rect 203616 88204 203668 88256
rect 87420 88136 87472 88188
rect 164884 88136 164936 88188
rect 110144 88068 110196 88120
rect 167828 88068 167880 88120
rect 135904 88000 135956 88052
rect 185676 88000 185728 88052
rect 121092 87932 121144 87984
rect 170496 87932 170548 87984
rect 300124 87660 300176 87712
rect 324320 87660 324372 87712
rect 3516 87592 3568 87644
rect 21364 87592 21416 87644
rect 185584 87592 185636 87644
rect 307300 87592 307352 87644
rect 63408 86912 63460 86964
rect 206376 86912 206428 86964
rect 274088 86912 274140 86964
rect 580172 86912 580224 86964
rect 99932 86844 99984 86896
rect 200764 86844 200816 86896
rect 117136 86776 117188 86828
rect 213276 86776 213328 86828
rect 102968 86708 103020 86760
rect 177396 86708 177448 86760
rect 122380 86640 122432 86692
rect 193864 86640 193916 86692
rect 252560 86232 252612 86284
rect 291936 86232 291988 86284
rect 67640 85484 67692 85536
rect 214840 85484 214892 85536
rect 85028 85416 85080 85468
rect 173440 85416 173492 85468
rect 96528 85348 96580 85400
rect 167920 85348 167972 85400
rect 118240 85280 118292 85332
rect 188436 85280 188488 85332
rect 135076 85212 135128 85264
rect 203524 85212 203576 85264
rect 116768 85144 116820 85196
rect 169116 85144 169168 85196
rect 238760 84872 238812 84924
rect 295432 84872 295484 84924
rect 179236 84804 179288 84856
rect 267832 84804 267884 84856
rect 64696 84124 64748 84176
rect 193956 84124 194008 84176
rect 112444 84056 112496 84108
rect 214656 84056 214708 84108
rect 119988 83988 120040 84040
rect 210516 83988 210568 84040
rect 106188 83920 106240 83972
rect 173256 83920 173308 83972
rect 129648 83852 129700 83904
rect 167644 83852 167696 83904
rect 285772 83512 285824 83564
rect 293040 83512 293092 83564
rect 176476 83444 176528 83496
rect 313280 83444 313332 83496
rect 100668 82764 100720 82816
rect 189908 82764 189960 82816
rect 126888 82696 126940 82748
rect 209044 82696 209096 82748
rect 115756 82628 115808 82680
rect 196808 82628 196860 82680
rect 86776 82560 86828 82612
rect 166540 82560 166592 82612
rect 103428 82492 103480 82544
rect 171876 82492 171928 82544
rect 198096 82220 198148 82272
rect 260104 82220 260156 82272
rect 216036 82152 216088 82204
rect 327080 82152 327132 82204
rect 191104 82084 191156 82136
rect 323584 82084 323636 82136
rect 45192 81336 45244 81388
rect 322940 81336 322992 81388
rect 92388 81268 92440 81320
rect 192760 81268 192812 81320
rect 95056 81200 95108 81252
rect 188528 81200 188580 81252
rect 131028 81132 131080 81184
rect 211896 81132 211948 81184
rect 120816 81064 120868 81116
rect 187148 81064 187200 81116
rect 35808 79976 35860 80028
rect 321836 79976 321888 80028
rect 102048 79908 102100 79960
rect 188344 79908 188396 79960
rect 120724 79840 120776 79892
rect 205088 79840 205140 79892
rect 97816 79772 97868 79824
rect 178684 79772 178736 79824
rect 99104 79704 99156 79756
rect 171968 79704 172020 79756
rect 39856 78616 39908 78668
rect 318064 78616 318116 78668
rect 97908 78548 97960 78600
rect 189816 78548 189868 78600
rect 125508 78480 125560 78532
rect 211988 78480 212040 78532
rect 118608 78412 118660 78464
rect 192668 78412 192720 78464
rect 99288 77188 99340 77240
rect 184296 77188 184348 77240
rect 114468 77120 114520 77172
rect 169024 77120 169076 77172
rect 115940 76576 115992 76628
rect 301780 76576 301832 76628
rect 80060 76508 80112 76560
rect 304540 76508 304592 76560
rect 308404 76508 308456 76560
rect 316132 76508 316184 76560
rect 93768 75828 93820 75880
rect 174636 75828 174688 75880
rect 111708 75760 111760 75812
rect 185768 75760 185820 75812
rect 184940 75216 184992 75268
rect 315304 75216 315356 75268
rect 98000 75148 98052 75200
rect 285128 75148 285180 75200
rect 127624 74468 127676 74520
rect 207756 74468 207808 74520
rect 81440 73856 81492 73908
rect 305736 73856 305788 73908
rect 6920 73788 6972 73840
rect 293408 73788 293460 73840
rect 309876 73652 309928 73704
rect 317420 73652 317472 73704
rect 356704 73108 356756 73160
rect 580172 73108 580224 73160
rect 85580 72496 85632 72548
rect 279516 72496 279568 72548
rect 46940 72428 46992 72480
rect 296168 72428 296220 72480
rect 3424 71680 3476 71732
rect 43444 71680 43496 71732
rect 113180 71136 113232 71188
rect 297548 71136 297600 71188
rect 44180 71068 44232 71120
rect 261668 71068 261720 71120
rect 37280 71000 37332 71052
rect 304448 71000 304500 71052
rect 51080 69640 51132 69692
rect 294880 69640 294932 69692
rect 92480 68348 92532 68400
rect 294696 68348 294748 68400
rect 57980 68280 58032 68332
rect 303160 68280 303212 68332
rect 99380 66920 99432 66972
rect 278320 66920 278372 66972
rect 64880 66852 64932 66904
rect 296076 66852 296128 66904
rect 106280 65560 106332 65612
rect 267004 65560 267056 65612
rect 69020 65492 69072 65544
rect 305920 65492 305972 65544
rect 71780 64200 71832 64252
rect 261576 64200 261628 64252
rect 34520 64132 34572 64184
rect 297640 64132 297692 64184
rect 110420 62840 110472 62892
rect 250628 62840 250680 62892
rect 117320 62772 117372 62824
rect 290556 62772 290608 62824
rect 82820 61412 82872 61464
rect 267096 61412 267148 61464
rect 67640 61344 67692 61396
rect 301596 61344 301648 61396
rect 359464 60664 359516 60716
rect 580172 60664 580224 60716
rect 85672 59984 85724 60036
rect 303068 59984 303120 60036
rect 3056 59304 3108 59356
rect 58624 59304 58676 59356
rect 120080 58692 120132 58744
rect 272524 58692 272576 58744
rect 89720 58624 89772 58676
rect 300400 58624 300452 58676
rect 74540 57264 74592 57316
rect 282276 57264 282328 57316
rect 93860 57196 93912 57248
rect 305828 57196 305880 57248
rect 96620 55904 96672 55956
rect 271236 55904 271288 55956
rect 70400 55836 70452 55888
rect 280988 55836 281040 55888
rect 100760 54544 100812 54596
rect 299020 54544 299072 54596
rect 63500 54476 63552 54528
rect 283840 54476 283892 54528
rect 103520 53116 103572 53168
rect 304356 53116 304408 53168
rect 60740 53048 60792 53100
rect 285036 53048 285088 53100
rect 107660 51756 107712 51808
rect 275376 51756 275428 51808
rect 4160 51688 4212 51740
rect 307208 51688 307260 51740
rect 84200 50396 84252 50448
rect 298928 50396 298980 50448
rect 44272 50328 44324 50380
rect 262956 50328 263008 50380
rect 102140 49036 102192 49088
rect 250444 49036 250496 49088
rect 124220 48968 124272 49020
rect 280896 48968 280948 49020
rect 30380 47608 30432 47660
rect 268476 47608 268528 47660
rect 49700 47540 49752 47592
rect 307116 47540 307168 47592
rect 353944 46860 353996 46912
rect 580172 46860 580224 46912
rect 35992 46248 36044 46300
rect 287796 46248 287848 46300
rect 20720 46180 20772 46232
rect 289268 46180 289320 46232
rect 3424 45500 3476 45552
rect 18604 45500 18656 45552
rect 19340 44888 19392 44940
rect 260196 44888 260248 44940
rect 40040 44820 40092 44872
rect 294788 44820 294840 44872
rect 102232 43460 102284 43512
rect 287888 43460 287940 43512
rect 38660 43392 38712 43444
rect 269856 43392 269908 43444
rect 118700 42100 118752 42152
rect 300308 42100 300360 42152
rect 41420 42032 41472 42084
rect 282368 42032 282420 42084
rect 110512 40740 110564 40792
rect 304264 40740 304316 40792
rect 9680 40672 9732 40724
rect 289176 40672 289228 40724
rect 42800 39380 42852 39432
rect 278228 39380 278280 39432
rect 11060 39312 11112 39364
rect 274180 39312 274232 39364
rect 45560 37884 45612 37936
rect 273996 37884 274048 37936
rect 78680 36592 78732 36644
rect 301688 36592 301740 36644
rect 19432 36524 19484 36576
rect 271144 36524 271196 36576
rect 128360 35232 128412 35284
rect 216680 35232 216732 35284
rect 238024 35232 238076 35284
rect 251364 35232 251416 35284
rect 12440 35164 12492 35216
rect 294604 35164 294656 35216
rect 53840 33804 53892 33856
rect 293316 33804 293368 33856
rect 31760 33736 31812 33788
rect 286324 33736 286376 33788
rect 3516 33056 3568 33108
rect 46204 33056 46256 33108
rect 345664 33056 345716 33108
rect 579896 33056 579948 33108
rect 180800 32512 180852 32564
rect 261576 32512 261628 32564
rect 201500 32444 201552 32496
rect 343640 32444 343692 32496
rect 93952 32376 94004 32428
rect 300216 32376 300268 32428
rect 200120 31152 200172 31204
rect 311900 31152 311952 31204
rect 104900 31084 104952 31136
rect 290464 31084 290516 31136
rect 75920 31016 75972 31068
rect 276664 31016 276716 31068
rect 73160 29656 73212 29708
rect 269764 29656 269816 29708
rect 17960 29588 18012 29640
rect 284944 29588 284996 29640
rect 86960 28296 87012 28348
rect 261484 28296 261536 28348
rect 22100 28228 22152 28280
rect 307024 28228 307076 28280
rect 297364 27548 297416 27600
rect 299480 27548 299532 27600
rect 179328 26936 179380 26988
rect 273260 26936 273312 26988
rect 26240 26868 26292 26920
rect 250536 26868 250588 26920
rect 210424 25644 210476 25696
rect 324412 25644 324464 25696
rect 176568 25576 176620 25628
rect 296720 25576 296772 25628
rect 77300 25508 77352 25560
rect 273904 25508 273956 25560
rect 62120 24148 62172 24200
rect 302976 24148 303028 24200
rect 2872 24080 2924 24132
rect 262864 24080 262916 24132
rect 8300 22720 8352 22772
rect 298836 22720 298888 22772
rect 59360 21428 59412 21480
rect 292028 21428 292080 21480
rect 11152 21360 11204 21412
rect 253296 21360 253348 21412
rect 3424 20612 3476 20664
rect 32404 20612 32456 20664
rect 216128 20612 216180 20664
rect 579896 20612 579948 20664
rect 175188 20000 175240 20052
rect 262220 20000 262272 20052
rect 91100 19932 91152 19984
rect 283656 19932 283708 19984
rect 114560 18572 114612 18624
rect 283748 18572 283800 18624
rect 187700 17416 187752 17468
rect 253204 17416 253256 17468
rect 207020 17348 207072 17400
rect 345020 17348 345072 17400
rect 95240 17280 95292 17332
rect 302884 17280 302936 17332
rect 24860 17212 24912 17264
rect 256148 17212 256200 17264
rect 112352 15852 112404 15904
rect 305644 15852 305696 15904
rect 179420 14560 179472 14612
rect 306380 14560 306432 14612
rect 122288 14492 122340 14544
rect 256056 14492 256108 14544
rect 66720 14424 66772 14476
rect 293224 14424 293276 14476
rect 119896 13064 119948 13116
rect 264336 13064 264388 13116
rect 179512 11840 179564 11892
rect 294880 11840 294932 11892
rect 109040 11772 109092 11824
rect 265716 11772 265768 11824
rect 33600 11704 33652 11756
rect 292120 11704 292172 11756
rect 112 10956 164 11008
rect 1308 10956 1360 11008
rect 251180 10956 251232 11008
rect 177948 10344 178000 10396
rect 287336 10344 287388 10396
rect 78128 10276 78180 10328
rect 295984 10276 296036 10328
rect 232504 9052 232556 9104
rect 281908 9052 281960 9104
rect 196624 8984 196676 9036
rect 260656 8984 260708 9036
rect 15936 8916 15988 8968
rect 289084 8916 289136 8968
rect 192484 7692 192536 7744
rect 299664 7692 299716 7744
rect 62028 7624 62080 7676
rect 298744 7624 298796 7676
rect 24216 7556 24268 7608
rect 279424 7556 279476 7608
rect 3424 6808 3476 6860
rect 22744 6808 22796 6860
rect 260104 6400 260156 6452
rect 284300 6400 284352 6452
rect 206284 6332 206336 6384
rect 266544 6332 266596 6384
rect 198740 6264 198792 6316
rect 276020 6264 276072 6316
rect 31668 6196 31720 6248
rect 136456 6196 136508 6248
rect 198004 6196 198056 6248
rect 292580 6196 292632 6248
rect 70308 6128 70360 6180
rect 301504 6128 301556 6180
rect 305552 6128 305604 6180
rect 338120 6128 338172 6180
rect 193220 4904 193272 4956
rect 247592 4904 247644 4956
rect 249984 4904 250036 4956
rect 265624 4904 265676 4956
rect 175096 4836 175148 4888
rect 304356 4836 304408 4888
rect 48964 4768 49016 4820
rect 278136 4768 278188 4820
rect 336004 4156 336056 4208
rect 340972 4156 341024 4208
rect 261576 4088 261628 4140
rect 268844 4088 268896 4140
rect 315304 4088 315356 4140
rect 316224 4088 316276 4140
rect 211804 3748 211856 3800
rect 245200 3748 245252 3800
rect 204904 3680 204956 3732
rect 242900 3680 242952 3732
rect 264888 3680 264940 3732
rect 271236 3680 271288 3732
rect 204168 3612 204220 3664
rect 248788 3612 248840 3664
rect 253204 3612 253256 3664
rect 261760 3612 261812 3664
rect 268384 3612 268436 3664
rect 283104 3612 283156 3664
rect 6460 3544 6512 3596
rect 56600 3544 56652 3596
rect 102140 3544 102192 3596
rect 103336 3544 103388 3596
rect 123484 3544 123536 3596
rect 228364 3544 228416 3596
rect 244096 3544 244148 3596
rect 255964 3544 256016 3596
rect 259460 3544 259512 3596
rect 275284 3544 275336 3596
rect 278044 3544 278096 3596
rect 288992 3544 289044 3596
rect 289728 3544 289780 3596
rect 293684 3544 293736 3596
rect 323584 3544 323636 3596
rect 337476 3544 337528 3596
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 19340 3476 19392 3528
rect 20260 3476 20312 3528
rect 35900 3476 35952 3528
rect 36820 3476 36872 3528
rect 52460 3476 52512 3528
rect 53380 3476 53432 3528
rect 57244 3476 57296 3528
rect 185584 3476 185636 3528
rect 189724 3476 189776 3528
rect 240508 3476 240560 3528
rect 252376 3476 252428 3528
rect 270500 3476 270552 3528
rect 28908 3408 28960 3460
rect 214564 3408 214616 3460
rect 215944 3408 215996 3460
rect 254676 3408 254728 3460
rect 264152 3408 264204 3460
rect 280804 3476 280856 3528
rect 287704 3476 287756 3528
rect 291384 3476 291436 3528
rect 299480 3476 299532 3528
rect 300768 3476 300820 3528
rect 316132 3476 316184 3528
rect 317328 3476 317380 3528
rect 324412 3476 324464 3528
rect 325608 3476 325660 3528
rect 332600 3476 332652 3528
rect 333888 3476 333940 3528
rect 280712 3408 280764 3460
rect 282184 3408 282236 3460
rect 291844 3408 291896 3460
rect 298468 3408 298520 3460
rect 309784 3408 309836 3460
rect 322112 3408 322164 3460
rect 326804 3340 326856 3392
rect 340880 3476 340932 3528
rect 323308 3272 323360 3324
rect 342260 3272 342312 3324
rect 264244 3204 264296 3256
rect 270040 3204 270092 3256
rect 330392 3204 330444 3256
rect 331496 3204 331548 3256
rect 308496 3136 308548 3188
rect 315028 3136 315080 3188
rect 345664 3136 345716 3188
rect 349252 3136 349304 3188
rect 249708 3000 249760 3052
rect 255872 3000 255924 3052
rect 235816 2932 235868 2984
rect 238024 2932 238076 2984
rect 337384 2932 337436 2984
rect 338672 2932 338724 2984
rect 56048 2048 56100 2100
rect 297456 2048 297508 2100
<< obsm1 >>
rect 68800 95100 164756 174600
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702710 8156 703520
rect 8116 702704 8168 702710
rect 8116 702646 8168 702652
rect 24320 700398 24348 703520
rect 37188 702840 37240 702846
rect 37188 702782 37240 702788
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 594114 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618662 3556 619103
rect 3516 618656 3568 618662
rect 3516 618598 3568 618604
rect 7564 618656 7616 618662
rect 7564 618598 7616 618604
rect 3514 606112 3570 606121
rect 3514 606047 3516 606056
rect 3568 606047 3570 606056
rect 3516 606018 3568 606024
rect 3424 594108 3476 594114
rect 3424 594050 3476 594056
rect 5448 587988 5500 587994
rect 5448 587930 5500 587936
rect 2872 583772 2924 583778
rect 2872 583714 2924 583720
rect 2884 580009 2912 583714
rect 2870 580000 2926 580009
rect 2870 579935 2926 579944
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3148 554736 3200 554742
rect 3148 554678 3200 554684
rect 3160 553897 3188 554678
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 3698 527912 3754 527921
rect 3698 527847 3754 527856
rect 3712 527202 3740 527847
rect 3700 527196 3752 527202
rect 3700 527138 3752 527144
rect 4068 527196 4120 527202
rect 4068 527138 4120 527144
rect 3424 516112 3476 516118
rect 3424 516054 3476 516060
rect 3436 514865 3464 516054
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3424 463684 3476 463690
rect 3424 463626 3476 463632
rect 3436 462641 3464 463626
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422294 3464 423535
rect 3436 422266 3556 422294
rect 3424 411256 3476 411262
rect 3424 411198 3476 411204
rect 3436 410553 3464 411198
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3528 407114 3556 422266
rect 3516 407108 3568 407114
rect 3516 407050 3568 407056
rect 3976 398132 4028 398138
rect 3976 398074 4028 398080
rect 3988 397497 4016 398074
rect 3974 397488 4030 397497
rect 3974 397423 4030 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 345704 3384 345710
rect 3332 345646 3384 345652
rect 3344 345409 3372 345646
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 319122 3464 319223
rect 3424 319116 3476 319122
rect 3424 319058 3476 319064
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 2688 293276 2740 293282
rect 2688 293218 2740 293224
rect 1306 177304 1362 177313
rect 1306 177239 1362 177248
rect 1320 11014 1348 177239
rect 2700 16561 2728 293218
rect 2870 293176 2926 293185
rect 2870 293111 2926 293120
rect 2884 291446 2912 293111
rect 2872 291440 2924 291446
rect 2872 291382 2924 291388
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3436 267034 3464 267135
rect 3424 267028 3476 267034
rect 3424 266970 3476 266976
rect 4080 262886 4108 527138
rect 5460 398138 5488 587930
rect 7576 543046 7604 618598
rect 8944 606076 8996 606082
rect 8944 606018 8996 606024
rect 7564 543040 7616 543046
rect 7564 542982 7616 542988
rect 7840 407108 7892 407114
rect 7840 407050 7892 407056
rect 7852 405754 7880 407050
rect 7840 405748 7892 405754
rect 7840 405690 7892 405696
rect 8208 405748 8260 405754
rect 8208 405690 8260 405696
rect 5448 398132 5500 398138
rect 5448 398074 5500 398080
rect 8220 297498 8248 405690
rect 8956 404530 8984 606018
rect 35808 589348 35860 589354
rect 35808 589290 35860 589296
rect 35164 586968 35216 586974
rect 35164 586910 35216 586916
rect 34428 586900 34480 586906
rect 34428 586842 34480 586848
rect 31024 585268 31076 585274
rect 31024 585210 31076 585216
rect 14464 565888 14516 565894
rect 14464 565830 14516 565836
rect 13084 477556 13136 477562
rect 13084 477498 13136 477504
rect 8944 404524 8996 404530
rect 8944 404466 8996 404472
rect 8944 319116 8996 319122
rect 8944 319058 8996 319064
rect 8956 311846 8984 319058
rect 8944 311840 8996 311846
rect 8944 311782 8996 311788
rect 8208 297492 8260 297498
rect 8208 297434 8260 297440
rect 4804 294024 4856 294030
rect 4804 293966 4856 293972
rect 4068 262880 4120 262886
rect 4068 262822 4120 262828
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 253978 3464 254079
rect 3424 253972 3476 253978
rect 3424 253914 3476 253920
rect 2962 241088 3018 241097
rect 2962 241023 3018 241032
rect 2976 237386 3004 241023
rect 2964 237380 3016 237386
rect 2964 237322 3016 237328
rect 3424 224256 3476 224262
rect 3424 224198 3476 224204
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3436 201929 3464 224198
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 4816 164150 4844 293966
rect 8944 291440 8996 291446
rect 8944 291382 8996 291388
rect 8956 244254 8984 291382
rect 13096 267034 13124 477498
rect 14476 404258 14504 565830
rect 27528 564460 27580 564466
rect 27528 564402 27580 564408
rect 22744 474768 22796 474774
rect 22744 474710 22796 474716
rect 17224 460964 17276 460970
rect 17224 460906 17276 460912
rect 17236 449886 17264 460906
rect 17224 449880 17276 449886
rect 17224 449822 17276 449828
rect 22756 428466 22784 474710
rect 22744 428460 22796 428466
rect 22744 428402 22796 428408
rect 17224 416832 17276 416838
rect 17224 416774 17276 416780
rect 14464 404252 14516 404258
rect 14464 404194 14516 404200
rect 17236 358766 17264 416774
rect 25504 398132 25556 398138
rect 25504 398074 25556 398080
rect 17224 358760 17276 358766
rect 17224 358702 17276 358708
rect 14464 347064 14516 347070
rect 14464 347006 14516 347012
rect 14476 345710 14504 347006
rect 14464 345704 14516 345710
rect 14464 345646 14516 345652
rect 14476 313954 14504 345646
rect 14464 313948 14516 313954
rect 14464 313890 14516 313896
rect 17224 290488 17276 290494
rect 17224 290430 17276 290436
rect 13084 267028 13136 267034
rect 13084 266970 13136 266976
rect 8944 244248 8996 244254
rect 8944 244190 8996 244196
rect 13096 234462 13124 266970
rect 14464 257372 14516 257378
rect 14464 257314 14516 257320
rect 13084 234456 13136 234462
rect 13084 234398 13136 234404
rect 13084 175976 13136 175982
rect 13084 175918 13136 175924
rect 2780 164144 2832 164150
rect 2780 164086 2832 164092
rect 4804 164144 4856 164150
rect 4804 164086 4856 164092
rect 2792 162897 2820 164086
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 13096 111790 13124 175918
rect 14476 137970 14504 257314
rect 17236 150414 17264 290430
rect 22744 279472 22796 279478
rect 22744 279414 22796 279420
rect 18604 263628 18656 263634
rect 18604 263570 18656 263576
rect 18616 215286 18644 263570
rect 21364 253224 21416 253230
rect 21364 253166 21416 253172
rect 18604 215280 18656 215286
rect 18604 215222 18656 215228
rect 18604 189848 18656 189854
rect 18604 189790 18656 189796
rect 17224 150408 17276 150414
rect 17224 150350 17276 150356
rect 14464 137964 14516 137970
rect 14464 137906 14516 137912
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 13084 111784 13136 111790
rect 13084 111726 13136 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3516 87644 3568 87650
rect 3516 87586 3568 87592
rect 3528 84697 3556 87586
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 6920 73840 6972 73846
rect 6920 73782 6972 73788
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 4160 51740 4212 51746
rect 4160 51682 4212 51688
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2778 37904 2834 37913
rect 2778 37839 2834 37848
rect 2686 16552 2742 16561
rect 2686 16487 2742 16496
rect 2700 15337 2728 16487
rect 1398 15328 1454 15337
rect 1398 15263 1454 15272
rect 2686 15328 2742 15337
rect 2686 15263 2742 15272
rect 112 11008 164 11014
rect 112 10950 164 10956
rect 1308 11008 1360 11014
rect 1308 10950 1360 10956
rect 124 354 152 10950
rect 542 354 654 480
rect 124 326 654 354
rect 1412 354 1440 15263
rect 2792 6914 2820 37839
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 2872 24132 2924 24138
rect 2872 24074 2924 24080
rect 2884 16574 2912 24074
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 51682
rect 6932 16574 6960 73782
rect 16578 62792 16634 62801
rect 16578 62727 16634 62736
rect 13818 59936 13874 59945
rect 13818 59871 13874 59880
rect 9680 40724 9732 40730
rect 9680 40666 9732 40672
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8312 16574 8340 22714
rect 2884 16546 3648 16574
rect 4172 16546 5304 16574
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 2792 6886 2912 6914
rect 2884 480 2912 6886
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 542 -960 654 326
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5276 480 5304 16546
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6472 480 6500 3538
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 40666
rect 11060 39364 11112 39370
rect 11060 39306 11112 39312
rect 11072 3534 11100 39306
rect 12440 35216 12492 35222
rect 12440 35158 12492 35164
rect 11152 21412 11204 21418
rect 11152 21354 11204 21360
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 21354
rect 12452 16574 12480 35158
rect 13832 16574 13860 59871
rect 16592 16574 16620 62727
rect 18616 45558 18644 189790
rect 21376 87650 21404 253166
rect 21364 87644 21416 87650
rect 21364 87586 21416 87592
rect 20720 46232 20772 46238
rect 20720 46174 20772 46180
rect 18604 45552 18656 45558
rect 18604 45494 18656 45500
rect 19340 44940 19392 44946
rect 19340 44882 19392 44888
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 16592 16546 17080 16574
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 480 15976 8910
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 29582
rect 19352 3534 19380 44882
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19444 480 19472 36518
rect 20732 16574 20760 46174
rect 22100 28280 22152 28286
rect 22100 28222 22152 28228
rect 22112 16574 22140 28222
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20272 354 20300 3470
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20272 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 22756 6866 22784 279414
rect 25516 239086 25544 398074
rect 26884 253972 26936 253978
rect 26884 253914 26936 253920
rect 25504 239080 25556 239086
rect 25504 239022 25556 239028
rect 26896 235890 26924 253914
rect 26884 235884 26936 235890
rect 26884 235826 26936 235832
rect 27540 232966 27568 564402
rect 31036 554742 31064 585210
rect 31666 558240 31722 558249
rect 31666 558175 31722 558184
rect 31024 554736 31076 554742
rect 31024 554678 31076 554684
rect 31576 538280 31628 538286
rect 31576 538222 31628 538228
rect 31588 360330 31616 538222
rect 31576 360324 31628 360330
rect 31576 360266 31628 360272
rect 31588 316742 31616 360266
rect 31576 316736 31628 316742
rect 31576 316678 31628 316684
rect 27528 232960 27580 232966
rect 27528 232902 27580 232908
rect 25504 213240 25556 213246
rect 25504 213182 25556 213188
rect 25516 97986 25544 213182
rect 25504 97980 25556 97986
rect 25504 97922 25556 97928
rect 30380 47660 30432 47666
rect 30380 47602 30432 47608
rect 26240 26920 26292 26926
rect 26240 26862 26292 26868
rect 24860 17264 24912 17270
rect 24860 17206 24912 17212
rect 24872 16574 24900 17206
rect 24872 16546 25360 16574
rect 24216 7608 24268 7614
rect 24216 7550 24268 7556
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 24228 480 24256 7550
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 26862
rect 27618 18592 27674 18601
rect 27618 18527 27674 18536
rect 27632 16574 27660 18527
rect 30392 16574 30420 47602
rect 27632 16546 27752 16574
rect 30392 16546 30880 16574
rect 27724 480 27752 16546
rect 30102 13016 30158 13025
rect 30102 12951 30158 12960
rect 28908 3460 28960 3466
rect 28908 3402 28960 3408
rect 28920 480 28948 3402
rect 30116 480 30144 12951
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31680 6254 31708 558175
rect 33048 554804 33100 554810
rect 33048 554746 33100 554752
rect 32956 488572 33008 488578
rect 32956 488514 33008 488520
rect 32404 299532 32456 299538
rect 32404 299474 32456 299480
rect 31760 33788 31812 33794
rect 31760 33730 31812 33736
rect 31772 16574 31800 33730
rect 32416 20670 32444 299474
rect 32968 281586 32996 488514
rect 33060 308446 33088 554746
rect 33048 308440 33100 308446
rect 33048 308382 33100 308388
rect 32956 281580 33008 281586
rect 32956 281522 33008 281528
rect 34440 242894 34468 586842
rect 35176 347070 35204 586910
rect 35164 347064 35216 347070
rect 35164 347006 35216 347012
rect 35820 290494 35848 589290
rect 37096 467900 37148 467906
rect 37096 467842 37148 467848
rect 35808 290488 35860 290494
rect 35808 290430 35860 290436
rect 35808 289128 35860 289134
rect 35808 289070 35860 289076
rect 35716 281580 35768 281586
rect 35716 281522 35768 281528
rect 34428 242888 34480 242894
rect 34428 242830 34480 242836
rect 35728 211818 35756 281522
rect 35716 211812 35768 211818
rect 35716 211754 35768 211760
rect 35820 80034 35848 289070
rect 37108 231674 37136 467842
rect 37200 407794 37228 702782
rect 40052 596834 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 63408 702772 63460 702778
rect 63408 702714 63460 702720
rect 53748 702568 53800 702574
rect 53748 702510 53800 702516
rect 48964 700392 49016 700398
rect 48964 700334 49016 700340
rect 45468 700324 45520 700330
rect 45468 700266 45520 700272
rect 43444 656940 43496 656946
rect 43444 656882 43496 656888
rect 40040 596828 40092 596834
rect 40040 596770 40092 596776
rect 42616 590844 42668 590850
rect 42616 590786 42668 590792
rect 39672 588192 39724 588198
rect 39672 588134 39724 588140
rect 38568 514820 38620 514826
rect 38568 514762 38620 514768
rect 37188 407788 37240 407794
rect 37188 407730 37240 407736
rect 37200 301481 37228 407730
rect 37186 301472 37242 301481
rect 37186 301407 37242 301416
rect 37096 231668 37148 231674
rect 37096 231610 37148 231616
rect 38580 229022 38608 514762
rect 39684 396982 39712 588134
rect 41326 586392 41382 586401
rect 41326 586327 41382 586336
rect 41236 585404 41288 585410
rect 41236 585346 41288 585352
rect 39856 552084 39908 552090
rect 39856 552026 39908 552032
rect 39764 423700 39816 423706
rect 39764 423642 39816 423648
rect 39672 396976 39724 396982
rect 39672 396918 39724 396924
rect 39672 368552 39724 368558
rect 39672 368494 39724 368500
rect 39684 244254 39712 368494
rect 39672 244248 39724 244254
rect 39672 244190 39724 244196
rect 39776 230450 39804 423642
rect 39868 358057 39896 552026
rect 39948 543040 40000 543046
rect 39948 542982 40000 542988
rect 39960 542434 39988 542982
rect 39948 542428 40000 542434
rect 39948 542370 40000 542376
rect 39854 358048 39910 358057
rect 39854 357983 39910 357992
rect 39854 284336 39910 284345
rect 39854 284271 39910 284280
rect 39764 230444 39816 230450
rect 39764 230386 39816 230392
rect 38568 229016 38620 229022
rect 38568 228958 38620 228964
rect 35808 80028 35860 80034
rect 35808 79970 35860 79976
rect 39868 78674 39896 284271
rect 39960 274650 39988 542370
rect 41144 388476 41196 388482
rect 41144 388418 41196 388424
rect 39948 274644 40000 274650
rect 39948 274586 40000 274592
rect 41156 237182 41184 388418
rect 41248 309806 41276 585346
rect 41236 309800 41288 309806
rect 41236 309742 41288 309748
rect 41236 278792 41288 278798
rect 41236 278734 41288 278740
rect 41144 237176 41196 237182
rect 41144 237118 41196 237124
rect 41248 181490 41276 278734
rect 41340 255270 41368 586327
rect 42524 414044 42576 414050
rect 42524 413986 42576 413992
rect 41420 311840 41472 311846
rect 41420 311782 41472 311788
rect 41432 311166 41460 311782
rect 41420 311160 41472 311166
rect 41420 311102 41472 311108
rect 41328 255264 41380 255270
rect 41328 255206 41380 255212
rect 42536 238746 42564 413986
rect 42628 311166 42656 590786
rect 42708 589416 42760 589422
rect 42708 589358 42760 589364
rect 42616 311160 42668 311166
rect 42616 311102 42668 311108
rect 42720 240786 42748 589358
rect 43456 402830 43484 656882
rect 45284 592136 45336 592142
rect 45284 592078 45336 592084
rect 44088 590776 44140 590782
rect 44088 590718 44140 590724
rect 43996 485852 44048 485858
rect 43996 485794 44048 485800
rect 43444 402824 43496 402830
rect 43444 402766 43496 402772
rect 43904 372224 43956 372230
rect 43904 372166 43956 372172
rect 43916 371278 43944 372166
rect 43904 371272 43956 371278
rect 43904 371214 43956 371220
rect 43916 297430 43944 371214
rect 44008 308514 44036 485794
rect 44100 403753 44128 590718
rect 44824 585472 44876 585478
rect 44824 585414 44876 585420
rect 44086 403744 44142 403753
rect 44086 403679 44142 403688
rect 44088 391332 44140 391338
rect 44088 391274 44140 391280
rect 43996 308508 44048 308514
rect 43996 308450 44048 308456
rect 43904 297424 43956 297430
rect 43904 297366 43956 297372
rect 43444 295452 43496 295458
rect 43444 295394 43496 295400
rect 42708 240780 42760 240786
rect 42708 240722 42760 240728
rect 42524 238740 42576 238746
rect 42524 238682 42576 238688
rect 41236 181484 41288 181490
rect 41236 181426 41288 181432
rect 39856 78668 39908 78674
rect 39856 78610 39908 78616
rect 43456 71738 43484 295394
rect 43996 284368 44048 284374
rect 43996 284310 44048 284316
rect 44008 209778 44036 284310
rect 44100 233034 44128 391274
rect 44836 372230 44864 585414
rect 45296 396914 45324 592078
rect 45376 470620 45428 470626
rect 45376 470562 45428 470568
rect 45284 396908 45336 396914
rect 45284 396850 45336 396856
rect 45284 394052 45336 394058
rect 45284 393994 45336 394000
rect 44824 372224 44876 372230
rect 44824 372166 44876 372172
rect 45192 251252 45244 251258
rect 45192 251194 45244 251200
rect 44088 233028 44140 233034
rect 44088 232970 44140 232976
rect 43996 209772 44048 209778
rect 43996 209714 44048 209720
rect 45204 81394 45232 251194
rect 45296 233102 45324 393994
rect 45388 237250 45416 470562
rect 45480 387802 45508 700266
rect 46204 683188 46256 683194
rect 46204 683130 46256 683136
rect 46216 529922 46244 683130
rect 48976 607170 49004 700334
rect 48964 607164 49016 607170
rect 48964 607106 49016 607112
rect 52276 607164 52328 607170
rect 52276 607106 52328 607112
rect 52288 605878 52316 607106
rect 52276 605872 52328 605878
rect 52276 605814 52328 605820
rect 46848 592204 46900 592210
rect 46848 592146 46900 592152
rect 46756 590708 46808 590714
rect 46756 590650 46808 590656
rect 46204 529916 46256 529922
rect 46204 529858 46256 529864
rect 46204 527196 46256 527202
rect 46204 527138 46256 527144
rect 46216 402966 46244 527138
rect 46664 437504 46716 437510
rect 46664 437446 46716 437452
rect 46204 402960 46256 402966
rect 46204 402902 46256 402908
rect 45468 387796 45520 387802
rect 45468 387738 45520 387744
rect 45480 249762 45508 387738
rect 45468 249756 45520 249762
rect 45468 249698 45520 249704
rect 46676 237318 46704 437446
rect 46768 356114 46796 590650
rect 46756 356108 46808 356114
rect 46756 356050 46808 356056
rect 46768 305658 46796 356050
rect 46756 305652 46808 305658
rect 46756 305594 46808 305600
rect 46860 302938 46888 592146
rect 48136 592068 48188 592074
rect 48136 592010 48188 592016
rect 48044 495508 48096 495514
rect 48044 495450 48096 495456
rect 48056 363662 48084 495450
rect 48148 400926 48176 592010
rect 52184 589484 52236 589490
rect 52184 589426 52236 589432
rect 48964 587920 49016 587926
rect 48964 587862 49016 587868
rect 48228 561740 48280 561746
rect 48228 561682 48280 561688
rect 48136 400920 48188 400926
rect 48136 400862 48188 400868
rect 48136 393984 48188 393990
rect 48136 393926 48188 393932
rect 48044 363656 48096 363662
rect 48044 363598 48096 363604
rect 46848 302932 46900 302938
rect 46848 302874 46900 302880
rect 46848 293344 46900 293350
rect 46848 293286 46900 293292
rect 46756 267776 46808 267782
rect 46756 267718 46808 267724
rect 46664 237312 46716 237318
rect 46664 237254 46716 237260
rect 45376 237244 45428 237250
rect 45376 237186 45428 237192
rect 46768 235958 46796 267718
rect 46756 235952 46808 235958
rect 46756 235894 46808 235900
rect 46768 234666 46796 235894
rect 46860 235754 46888 293286
rect 48044 289876 48096 289882
rect 48044 289818 48096 289824
rect 46848 235748 46900 235754
rect 46848 235690 46900 235696
rect 46204 234660 46256 234666
rect 46204 234602 46256 234608
rect 46756 234660 46808 234666
rect 46756 234602 46808 234608
rect 45284 233096 45336 233102
rect 45284 233038 45336 233044
rect 45192 81388 45244 81394
rect 45192 81330 45244 81336
rect 43444 71732 43496 71738
rect 43444 71674 43496 71680
rect 44180 71120 44232 71126
rect 44180 71062 44232 71068
rect 37280 71052 37332 71058
rect 37280 70994 37332 71000
rect 34520 64184 34572 64190
rect 34520 64126 34572 64132
rect 32404 20664 32456 20670
rect 32404 20606 32456 20612
rect 31772 16546 31984 16574
rect 31668 6248 31720 6254
rect 31668 6190 31720 6196
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 11756 33652 11762
rect 33600 11698 33652 11704
rect 33612 480 33640 11698
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 64126
rect 35898 48920 35954 48929
rect 35898 48855 35954 48864
rect 35912 3534 35940 48855
rect 35992 46300 36044 46306
rect 35992 46242 36044 46248
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36004 480 36032 46242
rect 37292 16574 37320 70994
rect 40040 44872 40092 44878
rect 40040 44814 40092 44820
rect 38660 43444 38712 43450
rect 38660 43386 38712 43392
rect 38672 16574 38700 43386
rect 40052 16574 40080 44814
rect 41420 42084 41472 42090
rect 41420 42026 41472 42032
rect 41432 16574 41460 42026
rect 42800 39432 42852 39438
rect 42800 39374 42852 39380
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36832 354 36860 3470
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 39374
rect 44192 6914 44220 71062
rect 44272 50380 44324 50386
rect 44272 50322 44324 50328
rect 44284 16574 44312 50322
rect 45560 37936 45612 37942
rect 45560 37878 45612 37884
rect 45572 16574 45600 37878
rect 46216 33114 46244 234602
rect 48056 205018 48084 289818
rect 48148 238950 48176 393926
rect 48240 249694 48268 561682
rect 48976 411262 49004 587862
rect 49516 586832 49568 586838
rect 49516 586774 49568 586780
rect 49424 428460 49476 428466
rect 49424 428402 49476 428408
rect 49436 427854 49464 428402
rect 49424 427848 49476 427854
rect 49424 427790 49476 427796
rect 48964 411256 49016 411262
rect 48964 411198 49016 411204
rect 49436 371890 49464 427790
rect 49424 371884 49476 371890
rect 49424 371826 49476 371832
rect 49424 352572 49476 352578
rect 49424 352514 49476 352520
rect 49436 266354 49464 352514
rect 49528 341465 49556 586774
rect 50344 585336 50396 585342
rect 50344 585278 50396 585284
rect 50986 585304 51042 585313
rect 49608 583840 49660 583846
rect 49608 583782 49660 583788
rect 49514 341456 49570 341465
rect 49514 341391 49570 341400
rect 49620 314022 49648 583782
rect 50356 463690 50384 585278
rect 50986 585239 51042 585248
rect 50436 501016 50488 501022
rect 50436 500958 50488 500964
rect 50344 463684 50396 463690
rect 50344 463626 50396 463632
rect 50448 404462 50476 500958
rect 50804 456816 50856 456822
rect 50804 456758 50856 456764
rect 50436 404456 50488 404462
rect 50436 404398 50488 404404
rect 49608 314016 49660 314022
rect 49608 313958 49660 313964
rect 50816 311234 50844 456758
rect 50896 441652 50948 441658
rect 50896 441594 50948 441600
rect 50804 311228 50856 311234
rect 50804 311170 50856 311176
rect 50908 295322 50936 441594
rect 51000 403850 51028 585239
rect 52092 460964 52144 460970
rect 52092 460906 52144 460912
rect 50988 403844 51040 403850
rect 50988 403786 51040 403792
rect 52104 366450 52132 460906
rect 52196 395350 52224 589426
rect 52288 399566 52316 605814
rect 53656 590912 53708 590918
rect 53656 590854 53708 590860
rect 53564 589620 53616 589626
rect 53564 589562 53616 589568
rect 52368 585200 52420 585206
rect 52368 585142 52420 585148
rect 52380 401713 52408 585142
rect 53472 529916 53524 529922
rect 53472 529858 53524 529864
rect 53484 528630 53512 529858
rect 53472 528624 53524 528630
rect 53472 528566 53524 528572
rect 52366 401704 52422 401713
rect 52366 401639 52422 401648
rect 52276 399560 52328 399566
rect 52276 399502 52328 399508
rect 52184 395344 52236 395350
rect 52184 395286 52236 395292
rect 52368 391264 52420 391270
rect 52368 391206 52420 391212
rect 52092 366444 52144 366450
rect 52092 366386 52144 366392
rect 52092 351212 52144 351218
rect 52092 351154 52144 351160
rect 50988 349852 51040 349858
rect 50988 349794 51040 349800
rect 50896 295316 50948 295322
rect 50896 295258 50948 295264
rect 49608 288448 49660 288454
rect 49608 288390 49660 288396
rect 49516 274712 49568 274718
rect 49516 274654 49568 274660
rect 49424 266348 49476 266354
rect 49424 266290 49476 266296
rect 48228 249688 48280 249694
rect 48228 249630 48280 249636
rect 48136 238944 48188 238950
rect 48136 238886 48188 238892
rect 48044 205012 48096 205018
rect 48044 204954 48096 204960
rect 49528 187066 49556 274654
rect 49620 192506 49648 288390
rect 50896 287088 50948 287094
rect 50896 287030 50948 287036
rect 50804 276072 50856 276078
rect 50804 276014 50856 276020
rect 50712 261520 50764 261526
rect 50712 261462 50764 261468
rect 50724 218754 50752 261462
rect 50712 218748 50764 218754
rect 50712 218690 50764 218696
rect 50816 214810 50844 276014
rect 50908 216102 50936 287030
rect 51000 247042 51028 349794
rect 52104 258058 52132 351154
rect 52184 277432 52236 277438
rect 52184 277374 52236 277380
rect 52092 258052 52144 258058
rect 52092 257994 52144 258000
rect 52104 257378 52132 257994
rect 52092 257372 52144 257378
rect 52092 257314 52144 257320
rect 50988 247036 51040 247042
rect 50988 246978 51040 246984
rect 50896 216096 50948 216102
rect 50896 216038 50948 216044
rect 50804 214804 50856 214810
rect 50804 214746 50856 214752
rect 52196 200841 52224 277374
rect 52276 260908 52328 260914
rect 52276 260850 52328 260856
rect 52288 218958 52316 260850
rect 52380 235822 52408 391206
rect 53484 366382 53512 528566
rect 53576 410038 53604 589562
rect 53564 410032 53616 410038
rect 53564 409974 53616 409980
rect 53562 405648 53618 405657
rect 53562 405583 53618 405592
rect 53576 400110 53604 405583
rect 53564 400104 53616 400110
rect 53564 400046 53616 400052
rect 53668 371958 53696 590854
rect 53760 465050 53788 702510
rect 63316 702500 63368 702506
rect 63316 702442 63368 702448
rect 55036 589688 55088 589694
rect 55036 589630 55088 589636
rect 54944 588056 54996 588062
rect 54944 587998 54996 588004
rect 53748 465044 53800 465050
rect 53748 464986 53800 464992
rect 53760 464953 53788 464986
rect 53746 464944 53802 464953
rect 53746 464879 53802 464888
rect 54852 444440 54904 444446
rect 54852 444382 54904 444388
rect 53748 410032 53800 410038
rect 53748 409974 53800 409980
rect 53760 405142 53788 409974
rect 53748 405136 53800 405142
rect 53748 405078 53800 405084
rect 53656 371952 53708 371958
rect 53656 371894 53708 371900
rect 53472 366376 53524 366382
rect 53472 366318 53524 366324
rect 54864 365090 54892 444382
rect 54956 403617 54984 587998
rect 55048 403782 55076 589630
rect 61936 589552 61988 589558
rect 61936 589494 61988 589500
rect 56416 588260 56468 588266
rect 56416 588202 56468 588208
rect 55128 568608 55180 568614
rect 55128 568550 55180 568556
rect 55036 403776 55088 403782
rect 55036 403718 55088 403724
rect 54942 403608 54998 403617
rect 54942 403543 54998 403552
rect 54852 365084 54904 365090
rect 54852 365026 54904 365032
rect 53748 365016 53800 365022
rect 53748 364958 53800 364964
rect 53564 298784 53616 298790
rect 53564 298726 53616 298732
rect 52460 290488 52512 290494
rect 52460 290430 52512 290436
rect 52472 289950 52500 290430
rect 52460 289944 52512 289950
rect 52460 289886 52512 289892
rect 53472 264988 53524 264994
rect 53472 264930 53524 264936
rect 52368 235816 52420 235822
rect 52368 235758 52420 235764
rect 52276 218952 52328 218958
rect 52276 218894 52328 218900
rect 53484 210458 53512 264930
rect 53576 241466 53604 298726
rect 53656 289944 53708 289950
rect 53656 289886 53708 289892
rect 53564 241460 53616 241466
rect 53564 241402 53616 241408
rect 53668 227730 53696 289886
rect 53760 280158 53788 364958
rect 55140 362234 55168 568550
rect 55864 501016 55916 501022
rect 55864 500958 55916 500964
rect 55128 362228 55180 362234
rect 55128 362170 55180 362176
rect 55128 356720 55180 356726
rect 55128 356662 55180 356668
rect 54852 285728 54904 285734
rect 54852 285670 54904 285676
rect 53838 284336 53894 284345
rect 53838 284271 53840 284280
rect 53892 284271 53894 284280
rect 53840 284242 53892 284248
rect 53748 280152 53800 280158
rect 53748 280094 53800 280100
rect 53748 262268 53800 262274
rect 53748 262210 53800 262216
rect 53656 227724 53708 227730
rect 53656 227666 53708 227672
rect 53472 210452 53524 210458
rect 53472 210394 53524 210400
rect 52182 200832 52238 200841
rect 52182 200767 52238 200776
rect 49608 192500 49660 192506
rect 49608 192442 49660 192448
rect 53760 191214 53788 262210
rect 54864 225593 54892 285670
rect 55036 280220 55088 280226
rect 55036 280162 55088 280168
rect 54942 271824 54998 271833
rect 54942 271759 54998 271768
rect 54956 269822 54984 271759
rect 54944 269816 54996 269822
rect 54944 269758 54996 269764
rect 54850 225584 54906 225593
rect 54850 225519 54906 225528
rect 54956 207670 54984 269758
rect 55048 217462 55076 280162
rect 55140 238678 55168 356662
rect 55876 260846 55904 500958
rect 56232 491360 56284 491366
rect 56232 491302 56284 491308
rect 55864 260840 55916 260846
rect 55864 260782 55916 260788
rect 56244 238785 56272 491302
rect 56428 405074 56456 588202
rect 60096 588124 60148 588130
rect 60096 588066 60148 588072
rect 60004 586764 60056 586770
rect 60004 586706 60056 586712
rect 58622 586664 58678 586673
rect 58622 586599 58678 586608
rect 57888 583908 57940 583914
rect 57888 583850 57940 583856
rect 57794 583808 57850 583817
rect 57704 583772 57756 583778
rect 57900 583778 57928 583850
rect 57794 583743 57850 583752
rect 57888 583772 57940 583778
rect 57704 583714 57756 583720
rect 57244 535492 57296 535498
rect 57244 535434 57296 535440
rect 56416 405068 56468 405074
rect 56416 405010 56468 405016
rect 57256 278798 57284 535434
rect 57716 433294 57744 583714
rect 57704 433288 57756 433294
rect 57704 433230 57756 433236
rect 57808 412634 57836 583743
rect 57888 583714 57940 583720
rect 57888 548412 57940 548418
rect 57888 548354 57940 548360
rect 57716 412606 57836 412634
rect 57336 405748 57388 405754
rect 57336 405690 57388 405696
rect 57348 402898 57376 405690
rect 57716 405006 57744 412606
rect 57704 405000 57756 405006
rect 57704 404942 57756 404948
rect 57336 402892 57388 402898
rect 57336 402834 57388 402840
rect 57244 278792 57296 278798
rect 57244 278734 57296 278740
rect 57796 271924 57848 271930
rect 57796 271866 57848 271872
rect 56324 270564 56376 270570
rect 56324 270506 56376 270512
rect 56230 238776 56286 238785
rect 56230 238711 56286 238720
rect 55128 238672 55180 238678
rect 55128 238614 55180 238620
rect 56336 234598 56364 270506
rect 57704 258188 57756 258194
rect 57704 258130 57756 258136
rect 56416 258120 56468 258126
rect 56416 258062 56468 258068
rect 56324 234592 56376 234598
rect 56324 234534 56376 234540
rect 55036 217456 55088 217462
rect 55036 217398 55088 217404
rect 54944 207664 54996 207670
rect 54944 207606 54996 207612
rect 56428 196654 56456 258062
rect 57716 202337 57744 258130
rect 57808 214674 57836 271866
rect 57900 238066 57928 548354
rect 58636 469849 58664 586599
rect 58716 583772 58768 583778
rect 58716 583714 58768 583720
rect 58728 516118 58756 583714
rect 59176 521688 59228 521694
rect 59176 521630 59228 521636
rect 58716 516112 58768 516118
rect 58716 516054 58768 516060
rect 58716 513936 58768 513942
rect 58716 513878 58768 513884
rect 58622 469840 58678 469849
rect 58622 469775 58678 469784
rect 58728 434625 58756 513878
rect 59084 481704 59136 481710
rect 59084 481646 59136 481652
rect 58714 434616 58770 434625
rect 58714 434551 58770 434560
rect 58992 417444 59044 417450
rect 58992 417386 59044 417392
rect 59004 355366 59032 417386
rect 59096 396778 59124 481646
rect 59084 396772 59136 396778
rect 59084 396714 59136 396720
rect 59188 373318 59216 521630
rect 59268 434784 59320 434790
rect 59268 434726 59320 434732
rect 59176 373312 59228 373318
rect 59176 373254 59228 373260
rect 58992 355360 59044 355366
rect 58992 355302 59044 355308
rect 59174 314800 59230 314809
rect 59174 314735 59230 314744
rect 59084 302320 59136 302326
rect 59084 302262 59136 302268
rect 58624 292664 58676 292670
rect 58624 292606 58676 292612
rect 57888 238060 57940 238066
rect 57888 238002 57940 238008
rect 57796 214668 57848 214674
rect 57796 214610 57848 214616
rect 57702 202328 57758 202337
rect 57702 202263 57758 202272
rect 56416 196648 56468 196654
rect 56416 196590 56468 196596
rect 53748 191208 53800 191214
rect 53748 191150 53800 191156
rect 49516 187060 49568 187066
rect 49516 187002 49568 187008
rect 52552 178016 52604 178022
rect 52552 177958 52604 177964
rect 52564 177313 52592 177958
rect 52550 177304 52606 177313
rect 52550 177239 52606 177248
rect 46940 72480 46992 72486
rect 46940 72422 46992 72428
rect 46204 33108 46256 33114
rect 46204 33050 46256 33056
rect 46952 16574 46980 72422
rect 51080 69692 51132 69698
rect 51080 69634 51132 69640
rect 49700 47592 49752 47598
rect 49700 47534 49752 47540
rect 49712 16574 49740 47534
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 4820 49016 4826
rect 48964 4762 49016 4768
rect 48976 480 49004 4762
rect 50172 480 50200 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 69634
rect 57980 68332 58032 68338
rect 57980 68274 58032 68280
rect 52458 58576 52514 58585
rect 52458 58511 52514 58520
rect 52472 3534 52500 58511
rect 53840 33856 53892 33862
rect 53840 33798 53892 33804
rect 52550 26888 52606 26897
rect 52550 26823 52606 26832
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 26823
rect 53852 16574 53880 33798
rect 57992 16574 58020 68274
rect 58636 59362 58664 292606
rect 59096 280090 59124 302262
rect 59084 280084 59136 280090
rect 59084 280026 59136 280032
rect 59096 279478 59124 280026
rect 59084 279472 59136 279478
rect 59084 279414 59136 279420
rect 59084 263628 59136 263634
rect 59084 263570 59136 263576
rect 58716 249892 58768 249898
rect 58716 249834 58768 249840
rect 58728 249694 58756 249834
rect 58716 249688 58768 249694
rect 58716 249630 58768 249636
rect 58728 220250 58756 249630
rect 59096 238882 59124 263570
rect 59084 238876 59136 238882
rect 59084 238818 59136 238824
rect 59188 238610 59216 314735
rect 59280 256018 59308 434726
rect 60016 417450 60044 586706
rect 60108 513942 60136 588066
rect 61382 585168 61438 585177
rect 61382 585103 61438 585112
rect 60738 568984 60794 568993
rect 60738 568919 60794 568928
rect 60752 568614 60780 568919
rect 60740 568608 60792 568614
rect 60740 568550 60792 568556
rect 60738 565584 60794 565593
rect 60738 565519 60794 565528
rect 60752 564466 60780 565519
rect 60740 564460 60792 564466
rect 60740 564402 60792 564408
rect 60738 562184 60794 562193
rect 60738 562119 60794 562128
rect 60752 561746 60780 562119
rect 60740 561740 60792 561746
rect 60740 561682 60792 561688
rect 60738 555384 60794 555393
rect 60738 555319 60794 555328
rect 60752 554810 60780 555319
rect 60740 554804 60792 554810
rect 60740 554746 60792 554752
rect 60738 552664 60794 552673
rect 60738 552599 60794 552608
rect 60752 552090 60780 552599
rect 60740 552084 60792 552090
rect 60740 552026 60792 552032
rect 60738 549264 60794 549273
rect 60738 549199 60794 549208
rect 60752 548418 60780 549199
rect 60740 548412 60792 548418
rect 60740 548354 60792 548360
rect 60738 542464 60794 542473
rect 60738 542399 60740 542408
rect 60792 542399 60794 542408
rect 60740 542370 60792 542376
rect 60738 539064 60794 539073
rect 60738 538999 60794 539008
rect 60752 538286 60780 538999
rect 60740 538280 60792 538286
rect 60740 538222 60792 538228
rect 60738 535664 60794 535673
rect 60738 535599 60794 535608
rect 60752 535498 60780 535599
rect 60740 535492 60792 535498
rect 60740 535434 60792 535440
rect 60738 528864 60794 528873
rect 60738 528799 60794 528808
rect 60752 528630 60780 528799
rect 60740 528624 60792 528630
rect 60740 528566 60792 528572
rect 60370 518664 60426 518673
rect 60370 518599 60426 518608
rect 60096 513936 60148 513942
rect 60096 513878 60148 513884
rect 60004 417444 60056 417450
rect 60004 417386 60056 417392
rect 60384 403714 60412 518599
rect 60738 515264 60794 515273
rect 60738 515199 60794 515208
rect 60752 514826 60780 515199
rect 60740 514820 60792 514826
rect 60740 514762 60792 514768
rect 60554 505064 60610 505073
rect 60554 504999 60610 505008
rect 60464 416764 60516 416770
rect 60464 416706 60516 416712
rect 60372 403708 60424 403714
rect 60372 403650 60424 403656
rect 60476 298858 60504 416706
rect 60568 377466 60596 504999
rect 60738 502344 60794 502353
rect 60738 502279 60794 502288
rect 60752 501022 60780 502279
rect 60740 501016 60792 501022
rect 60740 500958 60792 500964
rect 60738 495544 60794 495553
rect 60738 495479 60740 495488
rect 60792 495479 60794 495488
rect 60740 495450 60792 495456
rect 60738 492144 60794 492153
rect 60738 492079 60794 492088
rect 60752 491366 60780 492079
rect 60740 491360 60792 491366
rect 60740 491302 60792 491308
rect 61396 489914 61424 585103
rect 61658 522064 61714 522073
rect 61658 521999 61714 522008
rect 61672 521694 61700 521999
rect 61660 521688 61712 521694
rect 61660 521630 61712 521636
rect 61948 510513 61976 589494
rect 62764 586696 62816 586702
rect 62764 586638 62816 586644
rect 62026 545864 62082 545873
rect 62026 545799 62082 545808
rect 61934 510504 61990 510513
rect 61934 510439 61990 510448
rect 61934 508464 61990 508473
rect 61934 508399 61990 508408
rect 61212 489886 61424 489914
rect 60738 488744 60794 488753
rect 60738 488679 60794 488688
rect 60752 488578 60780 488679
rect 60740 488572 60792 488578
rect 60740 488514 60792 488520
rect 61212 485858 61240 489886
rect 61842 485888 61898 485897
rect 61200 485852 61252 485858
rect 61842 485823 61898 485832
rect 61200 485794 61252 485800
rect 61212 485353 61240 485794
rect 61198 485344 61254 485353
rect 61198 485279 61254 485288
rect 61566 481944 61622 481953
rect 61566 481879 61622 481888
rect 61580 481710 61608 481879
rect 61568 481704 61620 481710
rect 61568 481646 61620 481652
rect 60738 478544 60794 478553
rect 60738 478479 60794 478488
rect 60752 477562 60780 478479
rect 60740 477556 60792 477562
rect 60740 477498 60792 477504
rect 61382 475144 61438 475153
rect 61382 475079 61438 475088
rect 60922 471744 60978 471753
rect 60922 471679 60978 471688
rect 60936 470626 60964 471679
rect 60924 470620 60976 470626
rect 60924 470562 60976 470568
rect 60738 468344 60794 468353
rect 60738 468279 60794 468288
rect 60752 467906 60780 468279
rect 60740 467900 60792 467906
rect 60740 467842 60792 467848
rect 60740 465044 60792 465050
rect 60740 464986 60792 464992
rect 60752 464953 60780 464986
rect 60738 464944 60794 464953
rect 60738 464879 60794 464888
rect 60738 461544 60794 461553
rect 60738 461479 60794 461488
rect 60752 460970 60780 461479
rect 60740 460964 60792 460970
rect 60740 460906 60792 460912
rect 60738 458144 60794 458153
rect 60738 458079 60794 458088
rect 60752 456822 60780 458079
rect 60740 456816 60792 456822
rect 60740 456758 60792 456764
rect 61396 455394 61424 475079
rect 61856 473249 61884 485823
rect 61842 473240 61898 473249
rect 61842 473175 61898 473184
rect 60648 455388 60700 455394
rect 60648 455330 60700 455336
rect 61384 455388 61436 455394
rect 61384 455330 61436 455336
rect 60556 377460 60608 377466
rect 60556 377402 60608 377408
rect 60464 298852 60516 298858
rect 60464 298794 60516 298800
rect 60004 294160 60056 294166
rect 60004 294102 60056 294108
rect 59268 256012 59320 256018
rect 59268 255954 59320 255960
rect 59176 238604 59228 238610
rect 59176 238546 59228 238552
rect 58716 220244 58768 220250
rect 58716 220186 58768 220192
rect 60016 189038 60044 294102
rect 60556 255332 60608 255338
rect 60556 255274 60608 255280
rect 60464 241528 60516 241534
rect 60464 241470 60516 241476
rect 60476 227118 60504 241470
rect 60568 235278 60596 255274
rect 60660 238202 60688 455330
rect 61750 454744 61806 454753
rect 61750 454679 61806 454688
rect 60738 445224 60794 445233
rect 60738 445159 60794 445168
rect 60752 444446 60780 445159
rect 60740 444440 60792 444446
rect 60740 444382 60792 444388
rect 60738 441824 60794 441833
rect 60738 441759 60794 441768
rect 60752 441658 60780 441759
rect 60740 441652 60792 441658
rect 60740 441594 60792 441600
rect 60922 438424 60978 438433
rect 60922 438359 60978 438368
rect 60936 437510 60964 438359
rect 60924 437504 60976 437510
rect 60924 437446 60976 437452
rect 61566 435024 61622 435033
rect 61566 434959 61622 434968
rect 61580 434790 61608 434959
rect 61568 434784 61620 434790
rect 61568 434726 61620 434732
rect 60738 428224 60794 428233
rect 60738 428159 60794 428168
rect 60752 427854 60780 428159
rect 60740 427848 60792 427854
rect 60740 427790 60792 427796
rect 60738 424824 60794 424833
rect 60738 424759 60794 424768
rect 60752 423706 60780 424759
rect 60740 423700 60792 423706
rect 60740 423642 60792 423648
rect 60738 414624 60794 414633
rect 60738 414559 60794 414568
rect 60752 414050 60780 414559
rect 60740 414044 60792 414050
rect 60740 413986 60792 413992
rect 60738 407824 60794 407833
rect 60738 407759 60740 407768
rect 60792 407759 60794 407768
rect 60740 407730 60792 407736
rect 61764 399498 61792 454679
rect 61842 452024 61898 452033
rect 61842 451959 61898 451968
rect 61752 399492 61804 399498
rect 61752 399434 61804 399440
rect 61856 359417 61884 451959
rect 61842 359408 61898 359417
rect 61842 359343 61898 359352
rect 61844 270632 61896 270638
rect 61844 270574 61896 270580
rect 61752 261588 61804 261594
rect 61752 261530 61804 261536
rect 61764 239465 61792 261530
rect 61750 239456 61806 239465
rect 61750 239391 61806 239400
rect 60648 238196 60700 238202
rect 60648 238138 60700 238144
rect 60556 235272 60608 235278
rect 60556 235214 60608 235220
rect 61856 233238 61884 270574
rect 61948 261594 61976 508399
rect 62040 276146 62068 545799
rect 62302 418024 62358 418033
rect 62302 417959 62358 417968
rect 62316 416838 62344 417959
rect 62304 416832 62356 416838
rect 62304 416774 62356 416780
rect 62776 416770 62804 586638
rect 63224 585812 63276 585818
rect 63224 585754 63276 585760
rect 63038 498944 63094 498953
rect 63038 498879 63094 498888
rect 62856 433288 62908 433294
rect 62856 433230 62908 433236
rect 62868 417450 62896 433230
rect 62856 417444 62908 417450
rect 62856 417386 62908 417392
rect 62764 416764 62816 416770
rect 62764 416706 62816 416712
rect 62120 363656 62172 363662
rect 62120 363598 62172 363604
rect 62132 362982 62160 363598
rect 62120 362976 62172 362982
rect 62120 362918 62172 362924
rect 62764 362976 62816 362982
rect 62764 362918 62816 362924
rect 62028 276140 62080 276146
rect 62028 276082 62080 276088
rect 62028 269136 62080 269142
rect 62028 269078 62080 269084
rect 61936 261588 61988 261594
rect 61936 261530 61988 261536
rect 61936 253972 61988 253978
rect 61936 253914 61988 253920
rect 61844 233232 61896 233238
rect 61844 233174 61896 233180
rect 61948 231810 61976 253914
rect 61936 231804 61988 231810
rect 61936 231746 61988 231752
rect 60464 227112 60516 227118
rect 60464 227054 60516 227060
rect 62040 211954 62068 269078
rect 62120 262880 62172 262886
rect 62120 262822 62172 262828
rect 62132 260778 62160 262822
rect 62212 262200 62264 262206
rect 62212 262142 62264 262148
rect 62224 261526 62252 262142
rect 62212 261520 62264 261526
rect 62212 261462 62264 261468
rect 62120 260772 62172 260778
rect 62120 260714 62172 260720
rect 62120 255264 62172 255270
rect 62120 255206 62172 255212
rect 62132 254590 62160 255206
rect 62120 254584 62172 254590
rect 62120 254526 62172 254532
rect 62776 253910 62804 362918
rect 63052 262206 63080 498879
rect 63236 449954 63264 585754
rect 63328 525473 63356 702442
rect 63314 525464 63370 525473
rect 63314 525399 63370 525408
rect 63314 449984 63370 449993
rect 63224 449948 63276 449954
rect 63314 449919 63370 449928
rect 63224 449890 63276 449896
rect 63328 431954 63356 449919
rect 63420 438433 63448 702714
rect 63500 698964 63552 698970
rect 63500 698906 63552 698912
rect 63512 471753 63540 698906
rect 71792 599622 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 600982 88380 702406
rect 105464 699718 105492 703520
rect 130384 702636 130436 702642
rect 130384 702578 130436 702584
rect 100024 699712 100076 699718
rect 100024 699654 100076 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 88340 600976 88392 600982
rect 88340 600918 88392 600924
rect 71780 599616 71832 599622
rect 71780 599558 71832 599564
rect 100036 592686 100064 699654
rect 90180 592680 90232 592686
rect 90180 592622 90232 592628
rect 100024 592680 100076 592686
rect 100024 592622 100076 592628
rect 86500 590912 86552 590918
rect 86500 590854 86552 590860
rect 80152 586968 80204 586974
rect 80152 586910 80204 586916
rect 77576 586900 77628 586906
rect 77576 586842 77628 586848
rect 63592 586560 63644 586566
rect 63592 586502 63644 586508
rect 63604 583914 63632 586502
rect 71136 585472 71188 585478
rect 71136 585414 71188 585420
rect 67916 585404 67968 585410
rect 67916 585346 67968 585352
rect 67928 584868 67956 585346
rect 71148 584868 71176 585414
rect 77588 584868 77616 586842
rect 79416 586628 79468 586634
rect 79416 586570 79468 586576
rect 79428 585818 79456 586570
rect 79416 585812 79468 585818
rect 79416 585754 79468 585760
rect 80164 584868 80192 586910
rect 83370 586664 83426 586673
rect 83370 586599 83426 586608
rect 83384 584868 83412 586599
rect 86512 584882 86540 590854
rect 90192 588266 90220 592622
rect 102600 592204 102652 592210
rect 102600 592146 102652 592152
rect 90180 588260 90232 588266
rect 90180 588202 90232 588208
rect 90192 584882 90220 588202
rect 96252 586832 96304 586838
rect 96252 586774 96304 586780
rect 86512 584854 86618 584882
rect 89838 584854 90220 584882
rect 96264 584868 96292 586774
rect 99378 586392 99434 586401
rect 99378 586327 99434 586336
rect 99392 584882 99420 586327
rect 102612 584882 102640 592146
rect 112260 590844 112312 590850
rect 112260 590786 112312 590792
rect 105912 588192 105964 588198
rect 105912 588134 105964 588140
rect 99392 584854 99498 584882
rect 102612 584854 102718 584882
rect 105924 584868 105952 588134
rect 109132 586764 109184 586770
rect 109132 586706 109184 586712
rect 109144 584868 109172 586706
rect 112272 584882 112300 590786
rect 130396 590306 130424 702578
rect 137848 700330 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 702846 202828 703520
rect 202788 702840 202840 702846
rect 202788 702782 202840 702788
rect 210424 702704 210476 702710
rect 210424 702646 210476 702652
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 134156 592136 134208 592142
rect 134156 592078 134208 592084
rect 130384 590300 130436 590306
rect 130384 590242 130436 590248
rect 130936 590300 130988 590306
rect 130936 590242 130988 590248
rect 118700 589688 118752 589694
rect 118700 589630 118752 589636
rect 115572 586696 115624 586702
rect 115572 586638 115624 586644
rect 112272 584854 112378 584882
rect 115584 584868 115612 586638
rect 118712 584882 118740 589630
rect 121920 589620 121972 589626
rect 121920 589562 121972 589568
rect 121932 584882 121960 589562
rect 130948 589558 130976 590242
rect 130936 589552 130988 589558
rect 130936 589494 130988 589500
rect 127808 588124 127860 588130
rect 127808 588066 127860 588072
rect 125232 585200 125284 585206
rect 125232 585142 125284 585148
rect 118712 584854 118818 584882
rect 121932 584854 122038 584882
rect 125244 584868 125272 585142
rect 127820 584868 127848 588066
rect 130948 584882 130976 589494
rect 134168 584882 134196 592078
rect 153212 591326 153240 702406
rect 169772 595474 169800 702406
rect 175372 630692 175424 630698
rect 175372 630634 175424 630640
rect 169760 595468 169812 595474
rect 169760 595410 169812 595416
rect 153476 592068 153528 592074
rect 153476 592010 153528 592016
rect 153200 591320 153252 591326
rect 153200 591262 153252 591268
rect 143816 590776 143868 590782
rect 143816 590718 143868 590724
rect 140596 589484 140648 589490
rect 140596 589426 140648 589432
rect 137468 586628 137520 586634
rect 137468 586570 137520 586576
rect 130948 584854 131054 584882
rect 134168 584854 134274 584882
rect 137480 584868 137508 586570
rect 140608 584882 140636 589426
rect 143828 584882 143856 590718
rect 147128 587988 147180 587994
rect 147128 587930 147180 587936
rect 140608 584854 140714 584882
rect 143828 584854 143934 584882
rect 147140 584868 147168 587930
rect 150348 586560 150400 586566
rect 150348 586502 150400 586508
rect 150360 584868 150388 586502
rect 153488 584882 153516 592010
rect 159916 590708 159968 590714
rect 159916 590650 159968 590656
rect 156696 589416 156748 589422
rect 156696 589358 156748 589364
rect 156708 584882 156736 589358
rect 159928 584882 159956 590650
rect 163136 589348 163188 589354
rect 163136 589290 163188 589296
rect 163148 584882 163176 589290
rect 172888 586560 172940 586566
rect 172888 586502 172940 586508
rect 169666 585440 169722 585449
rect 169666 585375 169722 585384
rect 166448 585200 166500 585206
rect 166448 585142 166500 585148
rect 153488 584854 153594 584882
rect 156708 584854 156814 584882
rect 159928 584854 160034 584882
rect 163148 584854 163254 584882
rect 166460 584868 166488 585142
rect 169680 584868 169708 585375
rect 172900 585342 172928 586502
rect 172888 585336 172940 585342
rect 172888 585278 172940 585284
rect 172900 584868 172928 585278
rect 175384 584882 175412 630634
rect 185032 605872 185084 605878
rect 185032 605814 185084 605820
rect 181904 586628 181956 586634
rect 181904 586570 181956 586576
rect 178682 585304 178738 585313
rect 178682 585239 178738 585248
rect 175384 584854 175490 584882
rect 178696 584868 178724 585239
rect 181916 584868 181944 586570
rect 185044 584882 185072 605814
rect 201408 589960 201460 589966
rect 201408 589902 201460 589908
rect 191564 588056 191616 588062
rect 191564 587998 191616 588004
rect 185044 584854 185150 584882
rect 191576 584868 191604 587998
rect 198004 587920 198056 587926
rect 198004 587862 198056 587868
rect 194784 585404 194836 585410
rect 194784 585346 194836 585352
rect 194796 584868 194824 585346
rect 198016 584868 198044 587862
rect 201420 586401 201448 589902
rect 210436 588062 210464 702646
rect 218992 698970 219020 703520
rect 235184 700330 235212 703520
rect 267660 702778 267688 703520
rect 267648 702772 267700 702778
rect 267648 702714 267700 702720
rect 248328 702704 248380 702710
rect 248328 702646 248380 702652
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 244280 700324 244332 700330
rect 244280 700266 244332 700272
rect 218980 698964 219032 698970
rect 218980 698906 219032 698912
rect 242808 683188 242860 683194
rect 242808 683130 242860 683136
rect 229744 632120 229796 632126
rect 229744 632062 229796 632068
rect 217324 596828 217376 596834
rect 217324 596770 217376 596776
rect 210424 588056 210476 588062
rect 210424 587998 210476 588004
rect 207664 586696 207716 586702
rect 207664 586638 207716 586644
rect 201406 586392 201462 586401
rect 201406 586327 201462 586336
rect 201420 584882 201448 586327
rect 201250 584854 201448 584882
rect 207676 584868 207704 586638
rect 210436 584882 210464 587998
rect 217336 586838 217364 596770
rect 220728 592680 220780 592686
rect 220728 592622 220780 592628
rect 217324 586832 217376 586838
rect 217324 586774 217376 586780
rect 214104 586764 214156 586770
rect 214104 586706 214156 586712
rect 210436 584854 210910 584882
rect 214116 584868 214144 586706
rect 217336 584868 217364 586774
rect 220740 585342 220768 592622
rect 229756 588198 229784 632062
rect 236644 600976 236696 600982
rect 236644 600918 236696 600924
rect 236656 589354 236684 600918
rect 236000 589348 236052 589354
rect 236000 589290 236052 589296
rect 236644 589348 236696 589354
rect 236644 589290 236696 589296
rect 229744 588192 229796 588198
rect 229744 588134 229796 588140
rect 226340 588124 226392 588130
rect 226340 588066 226392 588072
rect 220544 585336 220596 585342
rect 220544 585278 220596 585284
rect 220728 585336 220780 585342
rect 220728 585278 220780 585284
rect 220556 584868 220584 585278
rect 226352 584868 226380 588066
rect 229756 584882 229784 588134
rect 232778 586664 232834 586673
rect 232778 586599 232834 586608
rect 229586 584854 229784 584882
rect 232792 584868 232820 586599
rect 236012 584868 236040 589290
rect 242820 587994 242848 683130
rect 242808 587988 242860 587994
rect 242808 587930 242860 587936
rect 239220 586900 239272 586906
rect 239220 586842 239272 586848
rect 239232 584868 239260 586842
rect 242820 584882 242848 587930
rect 243176 586832 243228 586838
rect 243176 586774 243228 586780
rect 242992 586628 243044 586634
rect 242992 586570 243044 586576
rect 242466 584854 242848 584882
rect 64418 584624 64474 584633
rect 92754 584624 92810 584633
rect 64474 584582 64722 584610
rect 74000 584594 74382 584610
rect 73988 584588 74382 584594
rect 64418 584559 64474 584568
rect 74040 584582 74382 584588
rect 188066 584624 188122 584633
rect 92810 584582 93058 584610
rect 92754 584559 92810 584568
rect 223486 584624 223542 584633
rect 188122 584582 188370 584610
rect 204470 584594 204760 584610
rect 204470 584588 204772 584594
rect 204470 584582 204720 584588
rect 188066 584559 188122 584568
rect 73988 584530 74040 584536
rect 223146 584582 223486 584610
rect 223486 584559 223542 584568
rect 204720 584530 204772 584536
rect 63592 583908 63644 583914
rect 63592 583850 63644 583856
rect 243004 538214 243032 586570
rect 243188 581670 243216 586774
rect 243636 585404 243688 585410
rect 243636 585346 243688 585352
rect 243648 585177 243676 585346
rect 243266 585168 243322 585177
rect 243266 585103 243322 585112
rect 243634 585168 243690 585177
rect 243634 585103 243690 585112
rect 243176 581664 243228 581670
rect 243176 581606 243228 581612
rect 243280 578202 243308 585103
rect 243542 580952 243598 580961
rect 243542 580887 243598 580896
rect 243268 578196 243320 578202
rect 243268 578138 243320 578144
rect 243004 538186 243124 538214
rect 242912 532778 243032 532794
rect 242912 532772 243044 532778
rect 242912 532766 242992 532772
rect 63498 471744 63554 471753
rect 63498 471679 63554 471688
rect 63500 449948 63552 449954
rect 63500 449890 63552 449896
rect 63406 438424 63462 438433
rect 63406 438359 63462 438368
rect 63236 431926 63356 431954
rect 63236 429321 63264 431926
rect 63222 429312 63278 429321
rect 63512 429298 63540 449890
rect 63222 429247 63278 429256
rect 63420 429270 63540 429298
rect 63132 417444 63184 417450
rect 63132 417386 63184 417392
rect 63144 403646 63172 417386
rect 63224 416832 63276 416838
rect 63224 416774 63276 416780
rect 63132 403640 63184 403646
rect 63132 403582 63184 403588
rect 63236 396846 63264 416774
rect 63224 396840 63276 396846
rect 63224 396782 63276 396788
rect 63420 348430 63448 429270
rect 63682 410680 63738 410689
rect 63682 410615 63738 410624
rect 63500 404048 63552 404054
rect 63500 403990 63552 403996
rect 63408 348424 63460 348430
rect 63408 348366 63460 348372
rect 63316 262336 63368 262342
rect 63316 262278 63368 262284
rect 63040 262200 63092 262206
rect 63040 262142 63092 262148
rect 63132 254584 63184 254590
rect 63132 254526 63184 254532
rect 63144 254017 63172 254526
rect 63130 254008 63186 254017
rect 63130 253943 63186 253952
rect 62120 253904 62172 253910
rect 62120 253846 62172 253852
rect 62764 253904 62816 253910
rect 62764 253846 62816 253852
rect 62132 253230 62160 253846
rect 62120 253224 62172 253230
rect 62120 253166 62172 253172
rect 62120 251864 62172 251870
rect 62120 251806 62172 251812
rect 62132 251258 62160 251806
rect 62120 251252 62172 251258
rect 62120 251194 62172 251200
rect 63132 248464 63184 248470
rect 63132 248406 63184 248412
rect 62028 211948 62080 211954
rect 62028 211890 62080 211896
rect 63144 196722 63172 248406
rect 63224 247104 63276 247110
rect 63224 247046 63276 247052
rect 63236 229838 63264 247046
rect 63224 229832 63276 229838
rect 63224 229774 63276 229780
rect 63328 226302 63356 262278
rect 63406 252512 63462 252521
rect 63406 252447 63462 252456
rect 63420 251870 63448 252447
rect 63408 251864 63460 251870
rect 63408 251806 63460 251812
rect 63408 241596 63460 241602
rect 63408 241538 63460 241544
rect 63420 234530 63448 241538
rect 63512 239018 63540 403990
rect 63696 402974 63724 410615
rect 242806 405512 242862 405521
rect 242806 405447 242862 405456
rect 66904 405136 66956 405142
rect 63972 405062 64078 405090
rect 66272 405062 66654 405090
rect 236644 405136 236696 405142
rect 66904 405078 66956 405084
rect 63972 404054 64000 405062
rect 66166 404560 66222 404569
rect 66166 404495 66222 404504
rect 65522 404424 65578 404433
rect 66180 404394 66208 404495
rect 65522 404359 65578 404368
rect 66168 404388 66220 404394
rect 63960 404048 64012 404054
rect 63960 403990 64012 403996
rect 63696 402946 63908 402974
rect 63880 382974 63908 402946
rect 64144 396976 64196 396982
rect 64144 396918 64196 396924
rect 63868 382968 63920 382974
rect 63868 382910 63920 382916
rect 64156 294642 64184 396918
rect 64144 294636 64196 294642
rect 64144 294578 64196 294584
rect 64696 294636 64748 294642
rect 64696 294578 64748 294584
rect 64708 294545 64736 294578
rect 64694 294536 64750 294545
rect 64694 294471 64750 294480
rect 64604 276140 64656 276146
rect 64604 276082 64656 276088
rect 64616 242826 64644 276082
rect 65536 275534 65564 404359
rect 66168 404330 66220 404336
rect 66076 322244 66128 322250
rect 66076 322186 66128 322192
rect 65524 275528 65576 275534
rect 65524 275470 65576 275476
rect 65984 273284 66036 273290
rect 65984 273226 66036 273232
rect 64788 267844 64840 267850
rect 64788 267786 64840 267792
rect 64696 247172 64748 247178
rect 64696 247114 64748 247120
rect 64604 242820 64656 242826
rect 64604 242762 64656 242768
rect 63592 240780 63644 240786
rect 63592 240722 63644 240728
rect 63604 240174 63632 240722
rect 63592 240168 63644 240174
rect 63592 240110 63644 240116
rect 64604 240168 64656 240174
rect 64604 240110 64656 240116
rect 63500 239012 63552 239018
rect 63500 238954 63552 238960
rect 63408 234524 63460 234530
rect 63408 234466 63460 234472
rect 63316 226296 63368 226302
rect 63316 226238 63368 226244
rect 64616 221474 64644 240110
rect 64604 221468 64656 221474
rect 64604 221410 64656 221416
rect 63132 196716 63184 196722
rect 63132 196658 63184 196664
rect 60004 189032 60056 189038
rect 60004 188974 60056 188980
rect 64708 184414 64736 247114
rect 64696 184408 64748 184414
rect 64696 184350 64748 184356
rect 64800 180130 64828 267786
rect 65996 220114 66024 273226
rect 66088 246974 66116 322186
rect 66180 298178 66208 404330
rect 66168 298172 66220 298178
rect 66168 298114 66220 298120
rect 66180 284238 66208 298114
rect 66168 284232 66220 284238
rect 66168 284174 66220 284180
rect 66168 271992 66220 271998
rect 66168 271934 66220 271940
rect 66076 246968 66128 246974
rect 66076 246910 66128 246916
rect 66076 244316 66128 244322
rect 66076 244258 66128 244264
rect 65984 220108 66036 220114
rect 65984 220050 66036 220056
rect 66088 202230 66116 244258
rect 66180 206446 66208 271934
rect 66272 239970 66300 405062
rect 66260 239964 66312 239970
rect 66260 239906 66312 239912
rect 66916 238513 66944 405078
rect 69032 405062 69874 405090
rect 71976 405062 73094 405090
rect 75932 405062 76314 405090
rect 79336 405062 79534 405090
rect 80060 405068 80112 405074
rect 68284 403844 68336 403850
rect 68284 403786 68336 403792
rect 67638 399528 67694 399537
rect 67638 399463 67694 399472
rect 67652 306374 67680 399463
rect 67652 306346 67864 306374
rect 67546 296848 67602 296857
rect 67546 296783 67602 296792
rect 67456 291916 67508 291922
rect 67456 291858 67508 291864
rect 67468 288386 67496 291858
rect 67456 288380 67508 288386
rect 67456 288322 67508 288328
rect 67560 266665 67588 296783
rect 67730 291136 67786 291145
rect 67730 291071 67786 291080
rect 67638 290456 67694 290465
rect 67638 290391 67694 290400
rect 67652 289882 67680 290391
rect 67744 289950 67772 291071
rect 67732 289944 67784 289950
rect 67732 289886 67784 289892
rect 67640 289876 67692 289882
rect 67640 289818 67692 289824
rect 67730 289776 67786 289785
rect 67836 289762 67864 306346
rect 68296 305726 68324 403786
rect 68928 354816 68980 354822
rect 68928 354758 68980 354764
rect 68284 305720 68336 305726
rect 68284 305662 68336 305668
rect 68836 304292 68888 304298
rect 68836 304234 68888 304240
rect 68848 293146 68876 304234
rect 68836 293140 68888 293146
rect 68836 293082 68888 293088
rect 68940 293026 68968 354758
rect 69032 293350 69060 405062
rect 70584 366444 70636 366450
rect 70584 366386 70636 366392
rect 70596 365770 70624 366386
rect 70584 365764 70636 365770
rect 70584 365706 70636 365712
rect 70492 316736 70544 316742
rect 70492 316678 70544 316684
rect 69480 302932 69532 302938
rect 69480 302874 69532 302880
rect 69492 302258 69520 302874
rect 69112 302252 69164 302258
rect 69112 302194 69164 302200
rect 69480 302252 69532 302258
rect 69480 302194 69532 302200
rect 69020 293344 69072 293350
rect 69020 293286 69072 293292
rect 67786 289734 67864 289762
rect 68664 292998 68968 293026
rect 67730 289711 67786 289720
rect 67744 289134 67772 289711
rect 67732 289128 67784 289134
rect 67638 289096 67694 289105
rect 67732 289070 67784 289076
rect 67638 289031 67694 289040
rect 67652 288454 67680 289031
rect 67640 288448 67692 288454
rect 67640 288390 67692 288396
rect 67732 288380 67784 288386
rect 67732 288322 67784 288328
rect 67638 287736 67694 287745
rect 67638 287671 67694 287680
rect 67652 287094 67680 287671
rect 67640 287088 67692 287094
rect 67640 287030 67692 287036
rect 67744 286385 67772 288322
rect 67822 287056 67878 287065
rect 67822 286991 67878 287000
rect 67730 286376 67786 286385
rect 67730 286311 67786 286320
rect 67836 285734 67864 286991
rect 67824 285728 67876 285734
rect 67824 285670 67876 285676
rect 67640 284368 67692 284374
rect 67638 284336 67640 284345
rect 67692 284336 67694 284345
rect 67638 284271 67694 284280
rect 67732 284300 67784 284306
rect 67732 284242 67784 284248
rect 67640 284232 67692 284238
rect 67640 284174 67692 284180
rect 67652 282985 67680 284174
rect 67744 283665 67772 284242
rect 67730 283656 67786 283665
rect 67730 283591 67786 283600
rect 67638 282976 67694 282985
rect 67638 282911 67694 282920
rect 68664 281625 68692 292998
rect 68836 292936 68888 292942
rect 68742 292904 68798 292913
rect 68836 292878 68888 292884
rect 68742 292839 68798 292848
rect 68756 285025 68784 292839
rect 68742 285016 68798 285025
rect 68742 284951 68798 284960
rect 68650 281616 68706 281625
rect 68650 281551 68706 281560
rect 67640 281512 67692 281518
rect 67640 281454 67692 281460
rect 67652 280945 67680 281454
rect 67638 280936 67694 280945
rect 67638 280871 67694 280880
rect 67638 280256 67694 280265
rect 67638 280191 67640 280200
rect 67692 280191 67694 280200
rect 67640 280162 67692 280168
rect 67732 280152 67784 280158
rect 67732 280094 67784 280100
rect 67640 280084 67692 280090
rect 67640 280026 67692 280032
rect 67652 279585 67680 280026
rect 67638 279576 67694 279585
rect 67638 279511 67694 279520
rect 67744 278905 67772 280094
rect 67730 278896 67786 278905
rect 67730 278831 67786 278840
rect 67640 278724 67692 278730
rect 67640 278666 67692 278672
rect 67652 278225 67680 278666
rect 67638 278216 67694 278225
rect 67638 278151 67694 278160
rect 67638 277536 67694 277545
rect 67638 277471 67694 277480
rect 67652 277438 67680 277471
rect 67640 277432 67692 277438
rect 68848 277394 68876 292878
rect 69124 285705 69152 302194
rect 69204 292596 69256 292602
rect 69204 292538 69256 292544
rect 69110 285696 69166 285705
rect 69110 285631 69166 285640
rect 67640 277374 67692 277380
rect 68664 277366 68876 277394
rect 67730 276856 67786 276865
rect 67730 276791 67786 276800
rect 67638 276176 67694 276185
rect 67638 276111 67640 276120
rect 67692 276111 67694 276120
rect 67640 276082 67692 276088
rect 67744 276078 67772 276791
rect 67732 276072 67784 276078
rect 67732 276014 67784 276020
rect 68192 275528 68244 275534
rect 68190 275496 68192 275505
rect 68244 275496 68246 275505
rect 68190 275431 68246 275440
rect 67638 274816 67694 274825
rect 67638 274751 67694 274760
rect 67652 274718 67680 274751
rect 67640 274712 67692 274718
rect 67640 274654 67692 274660
rect 68008 274644 68060 274650
rect 68008 274586 68060 274592
rect 68020 274145 68048 274586
rect 68006 274136 68062 274145
rect 68006 274071 68062 274080
rect 67822 273456 67878 273465
rect 67822 273391 67878 273400
rect 67836 273290 67864 273391
rect 67824 273284 67876 273290
rect 67824 273226 67876 273232
rect 67638 272776 67694 272785
rect 67638 272711 67694 272720
rect 67652 271930 67680 272711
rect 67822 272096 67878 272105
rect 67822 272031 67878 272040
rect 67836 271998 67864 272031
rect 67824 271992 67876 271998
rect 67824 271934 67876 271940
rect 67640 271924 67692 271930
rect 67640 271866 67692 271872
rect 67730 271416 67786 271425
rect 67730 271351 67786 271360
rect 67638 270736 67694 270745
rect 67638 270671 67694 270680
rect 67652 270638 67680 270671
rect 67640 270632 67692 270638
rect 67640 270574 67692 270580
rect 67744 270570 67772 271351
rect 67732 270564 67784 270570
rect 67732 270506 67784 270512
rect 67730 270056 67786 270065
rect 67730 269991 67786 270000
rect 67640 269816 67692 269822
rect 67640 269758 67692 269764
rect 67652 269385 67680 269758
rect 67638 269376 67694 269385
rect 67638 269311 67694 269320
rect 67744 269142 67772 269991
rect 67732 269136 67784 269142
rect 67732 269078 67784 269084
rect 67730 268696 67786 268705
rect 67730 268631 67786 268640
rect 67638 268016 67694 268025
rect 67638 267951 67694 267960
rect 67652 267782 67680 267951
rect 67744 267850 67772 268631
rect 67732 267844 67784 267850
rect 67732 267786 67784 267792
rect 67640 267776 67692 267782
rect 67640 267718 67692 267724
rect 68664 267345 68692 277366
rect 68926 275496 68982 275505
rect 68926 275431 68982 275440
rect 68650 267336 68706 267345
rect 68650 267271 68706 267280
rect 67546 266656 67602 266665
rect 67546 266591 67602 266600
rect 67640 266348 67692 266354
rect 67640 266290 67692 266296
rect 67652 265305 67680 266290
rect 68098 265976 68154 265985
rect 68098 265911 68154 265920
rect 67638 265296 67694 265305
rect 67638 265231 67694 265240
rect 68112 264994 68140 265911
rect 68100 264988 68152 264994
rect 68100 264930 68152 264936
rect 67638 264616 67694 264625
rect 67638 264551 67694 264560
rect 67652 263634 67680 264551
rect 68834 263936 68890 263945
rect 68834 263871 68890 263880
rect 67640 263628 67692 263634
rect 67640 263570 67692 263576
rect 67730 263256 67786 263265
rect 67730 263191 67786 263200
rect 67638 262576 67694 262585
rect 67638 262511 67694 262520
rect 67652 262274 67680 262511
rect 67744 262342 67772 263191
rect 67732 262336 67784 262342
rect 67732 262278 67784 262284
rect 67640 262268 67692 262274
rect 67640 262210 67692 262216
rect 67732 262200 67784 262206
rect 67732 262142 67784 262148
rect 67638 261896 67694 261905
rect 67638 261831 67694 261840
rect 67652 261594 67680 261831
rect 67640 261588 67692 261594
rect 67640 261530 67692 261536
rect 67744 261225 67772 262142
rect 67730 261216 67786 261225
rect 67730 261151 67786 261160
rect 67732 260840 67784 260846
rect 67732 260782 67784 260788
rect 67640 260772 67692 260778
rect 67640 260714 67692 260720
rect 67652 260545 67680 260714
rect 67638 260536 67694 260545
rect 67638 260471 67694 260480
rect 67744 259865 67772 260782
rect 67730 259856 67786 259865
rect 67730 259791 67786 259800
rect 67730 259176 67786 259185
rect 67730 259111 67786 259120
rect 67638 258496 67694 258505
rect 67638 258431 67694 258440
rect 67652 258194 67680 258431
rect 67640 258188 67692 258194
rect 67640 258130 67692 258136
rect 67744 258126 67772 259111
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 67640 258052 67692 258058
rect 67640 257994 67692 258000
rect 67652 257825 67680 257994
rect 67638 257816 67694 257825
rect 67638 257751 67694 257760
rect 67638 256456 67694 256465
rect 67638 256391 67694 256400
rect 67652 255338 67680 256391
rect 67916 256012 67968 256018
rect 67916 255954 67968 255960
rect 67928 255785 67956 255954
rect 67914 255776 67970 255785
rect 67914 255711 67970 255720
rect 68742 255776 68798 255785
rect 68742 255711 68798 255720
rect 67640 255332 67692 255338
rect 67640 255274 67692 255280
rect 67730 255096 67786 255105
rect 67730 255031 67786 255040
rect 67640 254584 67692 254590
rect 67640 254526 67692 254532
rect 67652 254425 67680 254526
rect 67638 254416 67694 254425
rect 67638 254351 67694 254360
rect 67744 253978 67772 255031
rect 67732 253972 67784 253978
rect 67732 253914 67784 253920
rect 67640 253904 67692 253910
rect 67640 253846 67692 253852
rect 67652 253745 67680 253846
rect 67638 253736 67694 253745
rect 67638 253671 67694 253680
rect 67640 251864 67692 251870
rect 67640 251806 67692 251812
rect 67652 251705 67680 251806
rect 67638 251696 67694 251705
rect 67638 251631 67694 251640
rect 67638 251016 67694 251025
rect 67638 250951 67694 250960
rect 67546 250336 67602 250345
rect 67546 250271 67602 250280
rect 66996 242820 67048 242826
rect 66996 242762 67048 242768
rect 66902 238504 66958 238513
rect 66902 238439 66958 238448
rect 66168 206440 66220 206446
rect 66168 206382 66220 206388
rect 66076 202224 66128 202230
rect 66076 202166 66128 202172
rect 67008 188358 67036 242762
rect 67560 217394 67588 250271
rect 67652 249898 67680 250951
rect 67640 249892 67692 249898
rect 67640 249834 67692 249840
rect 67640 249756 67692 249762
rect 67640 249698 67692 249704
rect 67652 249665 67680 249698
rect 67638 249656 67694 249665
rect 67638 249591 67694 249600
rect 67638 248976 67694 248985
rect 67638 248911 67694 248920
rect 67652 248470 67680 248911
rect 67640 248464 67692 248470
rect 67640 248406 67692 248412
rect 67730 248296 67786 248305
rect 67730 248231 67786 248240
rect 67638 247616 67694 247625
rect 67638 247551 67694 247560
rect 67652 247178 67680 247551
rect 67640 247172 67692 247178
rect 67640 247114 67692 247120
rect 67744 247110 67772 248231
rect 67732 247104 67784 247110
rect 67732 247046 67784 247052
rect 67640 247036 67692 247042
rect 67640 246978 67692 246984
rect 67652 246945 67680 246978
rect 68192 246968 68244 246974
rect 67638 246936 67694 246945
rect 68192 246910 68244 246916
rect 67638 246871 67694 246880
rect 68204 246265 68232 246910
rect 68190 246256 68246 246265
rect 68190 246191 68246 246200
rect 68190 244896 68246 244905
rect 68190 244831 68246 244840
rect 68204 244322 68232 244831
rect 68192 244316 68244 244322
rect 68192 244258 68244 244264
rect 67640 244248 67692 244254
rect 67640 244190 67692 244196
rect 67652 243545 67680 244190
rect 67638 243536 67694 243545
rect 67638 243471 67694 243480
rect 67638 242856 67694 242865
rect 67638 242791 67694 242800
rect 67652 241602 67680 242791
rect 67730 242176 67786 242185
rect 67730 242111 67786 242120
rect 67640 241596 67692 241602
rect 67640 241538 67692 241544
rect 67744 241534 67772 242111
rect 67732 241528 67784 241534
rect 67638 241496 67694 241505
rect 67732 241470 67784 241476
rect 67638 241431 67640 241440
rect 67692 241431 67694 241440
rect 67640 241402 67692 241408
rect 67638 240816 67694 240825
rect 67638 240751 67694 240760
rect 67652 240174 67680 240751
rect 67640 240168 67692 240174
rect 67640 240110 67692 240116
rect 68756 231130 68784 255711
rect 68744 231124 68796 231130
rect 68744 231066 68796 231072
rect 68848 223582 68876 263871
rect 68836 223576 68888 223582
rect 68836 223518 68888 223524
rect 67548 217388 67600 217394
rect 67548 217330 67600 217336
rect 66996 188352 67048 188358
rect 66996 188294 67048 188300
rect 68940 181393 68968 275431
rect 69110 274136 69166 274145
rect 69110 274071 69166 274080
rect 69124 228954 69152 274071
rect 69216 265985 69244 292538
rect 70504 292369 70532 316678
rect 70596 306374 70624 365706
rect 71872 314696 71924 314702
rect 71872 314638 71924 314644
rect 70596 306346 70992 306374
rect 70676 294636 70728 294642
rect 70676 294578 70728 294584
rect 70490 292360 70546 292369
rect 70490 292295 70546 292304
rect 70688 291924 70716 294578
rect 70964 291938 70992 306346
rect 71778 295352 71834 295361
rect 71778 295287 71780 295296
rect 71832 295287 71834 295296
rect 71780 295258 71832 295264
rect 71884 291938 71912 314638
rect 71976 292602 72004 405062
rect 73158 404968 73214 404977
rect 73158 404903 73214 404912
rect 73172 315994 73200 404903
rect 73804 403776 73856 403782
rect 73804 403718 73856 403724
rect 73160 315988 73212 315994
rect 73160 315930 73212 315936
rect 73172 314702 73200 315930
rect 73160 314696 73212 314702
rect 73160 314638 73212 314644
rect 73816 303618 73844 403718
rect 75184 396908 75236 396914
rect 75184 396850 75236 396856
rect 75196 306474 75224 396850
rect 75932 388482 75960 405062
rect 79336 402830 79364 405062
rect 80060 405010 80112 405016
rect 79324 402824 79376 402830
rect 79324 402766 79376 402772
rect 76010 398168 76066 398177
rect 76010 398103 76066 398112
rect 75920 388476 75972 388482
rect 75920 388418 75972 388424
rect 75920 340196 75972 340202
rect 75920 340138 75972 340144
rect 75184 306468 75236 306474
rect 75184 306410 75236 306416
rect 73804 303612 73856 303618
rect 73804 303554 73856 303560
rect 73710 301200 73766 301209
rect 73710 301135 73766 301144
rect 72608 297492 72660 297498
rect 72608 297434 72660 297440
rect 71964 292596 72016 292602
rect 71964 292538 72016 292544
rect 70964 291910 71346 291938
rect 71884 291910 71990 291938
rect 72620 291924 72648 297434
rect 73252 294636 73304 294642
rect 73252 294578 73304 294584
rect 73264 291924 73292 294578
rect 73724 291922 73752 301135
rect 73894 295216 73950 295225
rect 73894 295151 73950 295160
rect 73908 291924 73936 295151
rect 75196 294642 75224 306410
rect 75184 294636 75236 294642
rect 75184 294578 75236 294584
rect 74540 294568 74592 294574
rect 74540 294510 74592 294516
rect 75826 294536 75882 294545
rect 74552 291924 74580 294510
rect 75826 294471 75882 294480
rect 75184 292732 75236 292738
rect 75184 292674 75236 292680
rect 75196 291924 75224 292674
rect 75840 291924 75868 294471
rect 75932 292074 75960 340138
rect 76024 294545 76052 398103
rect 79336 384334 79364 402766
rect 79324 384328 79376 384334
rect 79324 384270 79376 384276
rect 80072 356726 80100 405010
rect 82084 400920 82136 400926
rect 82084 400862 82136 400868
rect 80060 356720 80112 356726
rect 80060 356662 80112 356668
rect 79324 318096 79376 318102
rect 79324 318038 79376 318044
rect 79232 299668 79284 299674
rect 79232 299610 79284 299616
rect 77392 299600 77444 299606
rect 77392 299542 77444 299548
rect 76010 294536 76066 294545
rect 76010 294471 76066 294480
rect 77116 294024 77168 294030
rect 77116 293966 77168 293972
rect 75932 292046 76144 292074
rect 76116 291938 76144 292046
rect 73712 291916 73764 291922
rect 76116 291910 76498 291938
rect 77128 291924 77156 293966
rect 77404 291938 77432 299542
rect 78402 294264 78458 294273
rect 78402 294199 78458 294208
rect 77404 291910 77786 291938
rect 78416 291924 78444 294199
rect 79048 294092 79100 294098
rect 79048 294034 79100 294040
rect 79060 291924 79088 294034
rect 79244 291938 79272 299610
rect 79336 294098 79364 318038
rect 82096 307426 82124 400862
rect 82740 400178 82768 405076
rect 85592 405062 85974 405090
rect 88352 405062 89194 405090
rect 91112 405062 92414 405090
rect 95252 405062 95634 405090
rect 98012 405062 98854 405090
rect 82728 400172 82780 400178
rect 82728 400114 82780 400120
rect 82740 323610 82768 400114
rect 84844 399560 84896 399566
rect 84844 399502 84896 399508
rect 83464 345704 83516 345710
rect 83464 345646 83516 345652
rect 82728 323604 82780 323610
rect 82728 323546 82780 323552
rect 81440 307420 81492 307426
rect 81440 307362 81492 307368
rect 82084 307420 82136 307426
rect 82084 307362 82136 307368
rect 81452 306406 81480 307362
rect 81440 306400 81492 306406
rect 81440 306342 81492 306348
rect 80060 305652 80112 305658
rect 80060 305594 80112 305600
rect 79324 294092 79376 294098
rect 79324 294034 79376 294040
rect 80072 291938 80100 305594
rect 80980 294092 81032 294098
rect 80980 294034 81032 294040
rect 79244 291910 79718 291938
rect 80072 291910 80362 291938
rect 80992 291924 81020 294034
rect 81452 291938 81480 306342
rect 82268 295384 82320 295390
rect 82268 295326 82320 295332
rect 81452 291910 81650 291938
rect 82280 291924 82308 295326
rect 83476 294030 83504 345646
rect 84200 299804 84252 299810
rect 84200 299746 84252 299752
rect 83556 298240 83608 298246
rect 83556 298182 83608 298188
rect 83464 294024 83516 294030
rect 83464 293966 83516 293972
rect 82938 291922 83320 291938
rect 83568 291924 83596 298182
rect 84212 291924 84240 299746
rect 84856 292602 84884 399502
rect 85592 394058 85620 405062
rect 86224 395344 86276 395350
rect 86224 395286 86276 395292
rect 85580 394052 85632 394058
rect 85580 393994 85632 394000
rect 86236 306374 86264 395286
rect 88352 391338 88380 405062
rect 90362 398032 90418 398041
rect 90362 397967 90418 397976
rect 88340 391332 88392 391338
rect 88340 391274 88392 391280
rect 88340 329112 88392 329118
rect 88340 329054 88392 329060
rect 86236 306346 86448 306374
rect 86420 305114 86448 306346
rect 86408 305108 86460 305114
rect 86408 305050 86460 305056
rect 86132 296744 86184 296750
rect 86132 296686 86184 296692
rect 85488 294024 85540 294030
rect 85488 293966 85540 293972
rect 84844 292596 84896 292602
rect 84844 292538 84896 292544
rect 84856 291924 84884 292538
rect 85500 291924 85528 293966
rect 86144 291924 86172 296686
rect 86420 291938 86448 305050
rect 88064 295588 88116 295594
rect 88064 295530 88116 295536
rect 87420 295520 87472 295526
rect 87420 295462 87472 295468
rect 82938 291916 83332 291922
rect 82938 291910 83280 291916
rect 73712 291858 73764 291864
rect 86420 291910 86802 291938
rect 87432 291924 87460 295462
rect 88076 291924 88104 295530
rect 88352 291938 88380 329054
rect 90376 305017 90404 397967
rect 91112 375358 91140 405062
rect 95148 398812 95200 398818
rect 95148 398754 95200 398760
rect 91100 375352 91152 375358
rect 91100 375294 91152 375300
rect 92388 375352 92440 375358
rect 92388 375294 92440 375300
rect 92400 374066 92428 375294
rect 92388 374060 92440 374066
rect 92388 374002 92440 374008
rect 90456 352640 90508 352646
rect 90456 352582 90508 352588
rect 89718 305008 89774 305017
rect 89718 304943 89774 304952
rect 90362 305008 90418 305017
rect 90362 304943 90418 304952
rect 88982 303648 89038 303657
rect 88982 303583 88984 303592
rect 89036 303583 89038 303592
rect 88984 303554 89036 303560
rect 88996 291938 89024 303554
rect 89732 291938 89760 304943
rect 89812 294228 89864 294234
rect 89812 294170 89864 294176
rect 89824 293282 89852 294170
rect 90468 294030 90496 352582
rect 92400 302938 92428 374002
rect 95056 338972 95108 338978
rect 95056 338914 95108 338920
rect 92388 302932 92440 302938
rect 92388 302874 92440 302880
rect 92848 302388 92900 302394
rect 92848 302330 92900 302336
rect 91100 301504 91152 301510
rect 91100 301446 91152 301452
rect 90640 296812 90692 296818
rect 90640 296754 90692 296760
rect 90456 294024 90508 294030
rect 90456 293966 90508 293972
rect 89812 293276 89864 293282
rect 89812 293218 89864 293224
rect 88352 291910 88734 291938
rect 88996 291910 89378 291938
rect 89732 291910 90022 291938
rect 90652 291924 90680 296754
rect 91112 291938 91140 301446
rect 91744 298376 91796 298382
rect 91744 298318 91796 298324
rect 91756 294574 91784 298318
rect 91744 294568 91796 294574
rect 91744 294510 91796 294516
rect 92480 294160 92532 294166
rect 92480 294102 92532 294108
rect 91928 294024 91980 294030
rect 91928 293966 91980 293972
rect 91112 291910 91310 291938
rect 91940 291924 91968 293966
rect 92492 292874 92520 294102
rect 92480 292868 92532 292874
rect 92480 292810 92532 292816
rect 92492 291938 92520 292810
rect 92860 291938 92888 302330
rect 94136 300620 94188 300626
rect 94136 300562 94188 300568
rect 93860 294160 93912 294166
rect 93860 294102 93912 294108
rect 92492 291910 92598 291938
rect 92860 291910 93242 291938
rect 93872 291924 93900 294102
rect 94148 291938 94176 300562
rect 95068 297498 95096 338914
rect 95160 300626 95188 398754
rect 95252 393990 95280 405062
rect 96528 404524 96580 404530
rect 96528 404466 96580 404472
rect 96540 398818 96568 404466
rect 96528 398812 96580 398818
rect 96528 398754 96580 398760
rect 95240 393984 95292 393990
rect 95240 393926 95292 393932
rect 98012 391270 98040 405062
rect 98736 403708 98788 403714
rect 98736 403650 98788 403656
rect 98644 396840 98696 396846
rect 98644 396782 98696 396788
rect 98000 391264 98052 391270
rect 98000 391206 98052 391212
rect 95882 380216 95938 380225
rect 95882 380151 95938 380160
rect 95148 300620 95200 300626
rect 95148 300562 95200 300568
rect 95160 299742 95188 300562
rect 95148 299736 95200 299742
rect 95148 299678 95200 299684
rect 95056 297492 95108 297498
rect 95056 297434 95108 297440
rect 95068 296714 95096 297434
rect 95068 296686 95188 296714
rect 94148 291910 94530 291938
rect 95160 291924 95188 296686
rect 95792 294636 95844 294642
rect 95792 294578 95844 294584
rect 95804 291924 95832 294578
rect 95896 294234 95924 380151
rect 96620 365084 96672 365090
rect 96620 365026 96672 365032
rect 96632 364478 96660 365026
rect 96620 364472 96672 364478
rect 96620 364414 96672 364420
rect 96632 306374 96660 364414
rect 98000 308168 98052 308174
rect 98000 308110 98052 308116
rect 98012 306374 98040 308110
rect 96632 306346 96752 306374
rect 98012 306346 98592 306374
rect 95884 294228 95936 294234
rect 95884 294170 95936 294176
rect 96436 294228 96488 294234
rect 96436 294170 96488 294176
rect 96448 291924 96476 294170
rect 96724 292670 96752 306346
rect 97264 305720 97316 305726
rect 97264 305662 97316 305668
rect 97276 300898 97304 305662
rect 97264 300892 97316 300898
rect 97264 300834 97316 300840
rect 96712 292664 96764 292670
rect 96712 292606 96764 292612
rect 96724 291938 96752 292606
rect 97276 291938 97304 300834
rect 98368 293276 98420 293282
rect 98368 293218 98420 293224
rect 98380 292670 98408 293218
rect 98368 292664 98420 292670
rect 98368 292606 98420 292612
rect 96724 291910 97106 291938
rect 97276 291910 97750 291938
rect 98380 291924 98408 292606
rect 98564 291938 98592 306346
rect 98656 293282 98684 396782
rect 98748 308174 98776 403650
rect 100668 402348 100720 402354
rect 100668 402290 100720 402296
rect 100680 318170 100708 402290
rect 102060 402286 102088 405076
rect 104164 405000 104216 405006
rect 104164 404942 104216 404948
rect 103518 403608 103574 403617
rect 103518 403543 103574 403552
rect 102048 402280 102100 402286
rect 102048 402222 102100 402228
rect 102784 401804 102836 401810
rect 102784 401746 102836 401752
rect 100760 362228 100812 362234
rect 100760 362170 100812 362176
rect 100772 361622 100800 362170
rect 100760 361616 100812 361622
rect 100760 361558 100812 361564
rect 100668 318164 100720 318170
rect 100668 318106 100720 318112
rect 98736 308168 98788 308174
rect 98736 308110 98788 308116
rect 98748 307834 98776 308110
rect 98736 307828 98788 307834
rect 98736 307770 98788 307776
rect 100772 295458 100800 361558
rect 102796 338978 102824 401746
rect 102784 338972 102836 338978
rect 102784 338914 102836 338920
rect 103532 303498 103560 403543
rect 103612 314084 103664 314090
rect 103612 314026 103664 314032
rect 103440 303470 103560 303498
rect 103440 296993 103468 303470
rect 103426 296984 103482 296993
rect 103426 296919 103482 296928
rect 102232 296880 102284 296886
rect 102232 296822 102284 296828
rect 100944 295656 100996 295662
rect 100944 295598 100996 295604
rect 100760 295452 100812 295458
rect 100760 295394 100812 295400
rect 98644 293276 98696 293282
rect 98644 293218 98696 293224
rect 99656 292800 99708 292806
rect 99656 292742 99708 292748
rect 98564 291910 99038 291938
rect 99668 291924 99696 292742
rect 100956 291924 100984 295598
rect 101588 295452 101640 295458
rect 101588 295394 101640 295400
rect 101600 291924 101628 295394
rect 102244 291924 102272 296822
rect 103518 295488 103574 295497
rect 103518 295423 103574 295432
rect 102902 291922 103192 291938
rect 103532 291924 103560 295423
rect 103624 293962 103652 314026
rect 104176 295497 104204 404942
rect 105280 404326 105308 405076
rect 105268 404320 105320 404326
rect 105268 404262 105320 404268
rect 105280 401810 105308 404262
rect 108500 402354 108528 405076
rect 108488 402348 108540 402354
rect 108488 402290 108540 402296
rect 105268 401804 105320 401810
rect 105268 401746 105320 401752
rect 111076 399566 111104 405076
rect 113192 405062 114310 405090
rect 111064 399560 111116 399566
rect 111064 399502 111116 399508
rect 108946 389872 109002 389881
rect 108946 389807 109002 389816
rect 105542 387016 105598 387025
rect 105542 386951 105598 386960
rect 104346 296984 104402 296993
rect 104346 296919 104402 296928
rect 104162 295488 104218 295497
rect 104162 295423 104218 295432
rect 103612 293956 103664 293962
rect 103612 293898 103664 293904
rect 104360 291938 104388 296919
rect 105452 294228 105504 294234
rect 105452 294170 105504 294176
rect 104532 293956 104584 293962
rect 104532 293898 104584 293904
rect 102902 291916 103204 291922
rect 102902 291910 103152 291916
rect 83280 291858 83332 291864
rect 104190 291910 104388 291938
rect 104544 291938 104572 293898
rect 104544 291910 104834 291938
rect 105464 291924 105492 294170
rect 105556 292777 105584 386951
rect 106280 323604 106332 323610
rect 106280 323546 106332 323552
rect 106292 321570 106320 323546
rect 106280 321564 106332 321570
rect 106280 321506 106332 321512
rect 106292 306374 106320 321506
rect 106292 306346 107056 306374
rect 106740 298308 106792 298314
rect 106740 298250 106792 298256
rect 105542 292768 105598 292777
rect 105542 292703 105598 292712
rect 106094 292768 106150 292777
rect 106094 292703 106150 292712
rect 106108 291924 106136 292703
rect 106752 291924 106780 298250
rect 107028 291938 107056 306346
rect 108960 300801 108988 389807
rect 113192 387802 113220 405062
rect 117516 402354 117544 405076
rect 120736 404530 120764 405076
rect 120724 404524 120776 404530
rect 120724 404466 120776 404472
rect 117504 402348 117556 402354
rect 117504 402290 117556 402296
rect 122104 402280 122156 402286
rect 122104 402222 122156 402228
rect 116584 401668 116636 401674
rect 116584 401610 116636 401616
rect 113180 387796 113232 387802
rect 113180 387738 113232 387744
rect 114468 387796 114520 387802
rect 114468 387738 114520 387744
rect 114480 387122 114508 387738
rect 114468 387116 114520 387122
rect 114468 387058 114520 387064
rect 109684 377460 109736 377466
rect 109684 377402 109736 377408
rect 109696 357202 109724 377402
rect 111708 376032 111760 376038
rect 111708 375974 111760 375980
rect 109040 357196 109092 357202
rect 109040 357138 109092 357144
rect 109684 357196 109736 357202
rect 109684 357138 109736 357144
rect 107658 300792 107714 300801
rect 107658 300727 107714 300736
rect 108946 300792 109002 300801
rect 108946 300727 109002 300736
rect 107672 291938 107700 300727
rect 108304 299872 108356 299878
rect 108304 299814 108356 299820
rect 108316 291938 108344 299814
rect 108960 299577 108988 300727
rect 108946 299568 109002 299577
rect 108946 299503 109002 299512
rect 109052 293962 109080 357138
rect 109696 356726 109724 357138
rect 109684 356720 109736 356726
rect 109684 356662 109736 356668
rect 110326 349752 110382 349761
rect 110326 349687 110382 349696
rect 110340 301073 110368 349687
rect 111720 301578 111748 375974
rect 113824 373312 113876 373318
rect 113824 373254 113876 373260
rect 112444 371952 112496 371958
rect 112444 371894 112496 371900
rect 111800 303000 111852 303006
rect 111800 302942 111852 302948
rect 110880 301572 110932 301578
rect 110880 301514 110932 301520
rect 111708 301572 111760 301578
rect 111708 301514 111760 301520
rect 109130 301064 109186 301073
rect 109130 300999 109186 301008
rect 110326 301064 110382 301073
rect 110326 300999 110382 301008
rect 109040 293956 109092 293962
rect 109040 293898 109092 293904
rect 109144 291938 109172 300999
rect 110604 295452 110656 295458
rect 110604 295394 110656 295400
rect 109684 293956 109736 293962
rect 109684 293898 109736 293904
rect 109696 291938 109724 293898
rect 107028 291910 107410 291938
rect 107672 291910 108054 291938
rect 108316 291910 108698 291938
rect 109144 291910 109342 291938
rect 109696 291910 109986 291938
rect 110616 291924 110644 295394
rect 110892 291938 110920 301514
rect 111812 299878 111840 302942
rect 111800 299872 111852 299878
rect 111800 299814 111852 299820
rect 112456 298897 112484 371894
rect 113178 354784 113234 354793
rect 113178 354719 113234 354728
rect 112442 298888 112498 298897
rect 112442 298823 112498 298832
rect 111890 294128 111946 294137
rect 111890 294063 111946 294072
rect 110892 291910 111274 291938
rect 111904 291924 111932 294063
rect 112562 291922 112852 291938
rect 113192 291924 113220 354719
rect 113836 306374 113864 373254
rect 113836 306346 114048 306374
rect 114020 303686 114048 306346
rect 114008 303680 114060 303686
rect 114008 303622 114060 303628
rect 113822 292632 113878 292641
rect 113822 292567 113878 292576
rect 113836 291924 113864 292567
rect 114020 291938 114048 303622
rect 115296 302932 115348 302938
rect 115296 302874 115348 302880
rect 115112 295724 115164 295730
rect 115112 295666 115164 295672
rect 112562 291916 112864 291922
rect 112562 291910 112812 291916
rect 103152 291858 103204 291864
rect 114020 291910 114494 291938
rect 115124 291924 115152 295666
rect 115308 291938 115336 302874
rect 116596 298110 116624 401610
rect 118606 400888 118662 400897
rect 118606 400823 118662 400832
rect 117964 356176 118016 356182
rect 117964 356118 118016 356124
rect 116676 311160 116728 311166
rect 116676 311102 116728 311108
rect 115940 298104 115992 298110
rect 115940 298046 115992 298052
rect 116584 298104 116636 298110
rect 116584 298046 116636 298052
rect 115952 294234 115980 298046
rect 115940 294228 115992 294234
rect 115940 294170 115992 294176
rect 116688 292942 116716 311102
rect 116768 309868 116820 309874
rect 116768 309810 116820 309816
rect 116780 295730 116808 309810
rect 117976 299538 118004 356118
rect 117964 299532 118016 299538
rect 117964 299474 118016 299480
rect 117976 296714 118004 299474
rect 117884 296686 118004 296714
rect 116768 295724 116820 295730
rect 116768 295666 116820 295672
rect 117686 295624 117742 295633
rect 117686 295559 117742 295568
rect 116676 292936 116728 292942
rect 116676 292878 116728 292884
rect 116688 291938 116716 292878
rect 115308 291910 115782 291938
rect 116426 291910 116716 291938
rect 117070 291922 117360 291938
rect 117700 291924 117728 295559
rect 117884 291938 117912 296686
rect 118620 295633 118648 400823
rect 120724 399492 120776 399498
rect 120724 399434 120776 399440
rect 118700 313948 118752 313954
rect 118700 313890 118752 313896
rect 118712 306374 118740 313890
rect 118712 306346 119200 306374
rect 118974 298888 119030 298897
rect 118974 298823 119030 298832
rect 118606 295624 118662 295633
rect 118606 295559 118662 295568
rect 117964 294092 118016 294098
rect 117964 294034 118016 294040
rect 117976 292097 118004 294034
rect 117962 292088 118018 292097
rect 117962 292023 118018 292032
rect 118988 291938 119016 298823
rect 119066 291952 119122 291961
rect 117070 291916 117372 291922
rect 117070 291910 117320 291916
rect 112812 291858 112864 291864
rect 117884 291910 118358 291938
rect 118988 291924 119066 291938
rect 119002 291910 119066 291924
rect 119172 291938 119200 306346
rect 120080 305040 120132 305046
rect 120080 304982 120132 304988
rect 119172 291910 119752 291938
rect 119066 291887 119122 291896
rect 117320 291858 117372 291864
rect 69308 291230 70058 291258
rect 69202 265976 69258 265985
rect 69202 265911 69258 265920
rect 69112 228948 69164 228954
rect 69112 228890 69164 228896
rect 69308 199510 69336 291230
rect 119724 267734 119752 291910
rect 120092 286385 120120 304982
rect 120172 298852 120224 298858
rect 120172 298794 120224 298800
rect 120078 286376 120134 286385
rect 120078 286311 120134 286320
rect 120184 280945 120212 298794
rect 120170 280936 120226 280945
rect 120170 280871 120226 280880
rect 119724 267706 119936 267734
rect 69662 243672 69718 243681
rect 69662 243607 69718 243616
rect 69676 242894 69704 243607
rect 69664 242888 69716 242894
rect 69664 242830 69716 242836
rect 69296 199504 69348 199510
rect 69296 199446 69348 199452
rect 69676 184278 69704 242830
rect 119908 242214 119936 267706
rect 120736 262274 120764 399434
rect 121460 384328 121512 384334
rect 121460 384270 121512 384276
rect 121472 383722 121500 384270
rect 121460 383716 121512 383722
rect 121460 383658 121512 383664
rect 121368 305652 121420 305658
rect 121368 305594 121420 305600
rect 121380 305046 121408 305594
rect 121368 305040 121420 305046
rect 121368 304982 121420 304988
rect 120816 291916 120868 291922
rect 120816 291858 120868 291864
rect 120724 262268 120776 262274
rect 120724 262210 120776 262216
rect 120724 253972 120776 253978
rect 120724 253914 120776 253920
rect 120632 251184 120684 251190
rect 120632 251126 120684 251132
rect 120644 251025 120672 251126
rect 120170 251016 120226 251025
rect 120170 250951 120226 250960
rect 120630 251016 120686 251025
rect 120630 250951 120686 250960
rect 119988 242276 120040 242282
rect 119988 242218 120040 242224
rect 119896 242208 119948 242214
rect 119896 242150 119948 242156
rect 119894 240952 119950 240961
rect 119894 240887 119950 240896
rect 70044 239018 70072 240108
rect 70688 239970 70716 240108
rect 70676 239964 70728 239970
rect 70676 239906 70728 239912
rect 70032 239012 70084 239018
rect 70032 238954 70084 238960
rect 70044 237454 70072 238954
rect 70032 237448 70084 237454
rect 70032 237390 70084 237396
rect 70688 219434 70716 239906
rect 71332 238134 71360 240108
rect 71320 238128 71372 238134
rect 71320 238070 71372 238076
rect 71044 237448 71096 237454
rect 71044 237390 71096 237396
rect 70412 219406 70716 219434
rect 70412 191146 70440 219406
rect 71056 217326 71084 237390
rect 71976 235754 72004 240108
rect 72620 238649 72648 240108
rect 72606 238640 72662 238649
rect 72606 238575 72662 238584
rect 72620 237153 72648 238575
rect 73068 238196 73120 238202
rect 73068 238138 73120 238144
rect 72606 237144 72662 237153
rect 72606 237079 72662 237088
rect 71964 235748 72016 235754
rect 71964 235690 72016 235696
rect 71976 234666 72004 235690
rect 71964 234660 72016 234666
rect 71964 234602 72016 234608
rect 72424 234660 72476 234666
rect 72424 234602 72476 234608
rect 71044 217320 71096 217326
rect 71044 217262 71096 217268
rect 72436 203590 72464 234602
rect 72424 203584 72476 203590
rect 72424 203526 72476 203532
rect 70400 191140 70452 191146
rect 70400 191082 70452 191088
rect 69664 184272 69716 184278
rect 69664 184214 69716 184220
rect 73080 182850 73108 238138
rect 73264 237182 73292 240108
rect 73908 238202 73936 240108
rect 74552 238785 74580 240108
rect 74538 238776 74594 238785
rect 75196 238754 75224 240108
rect 75840 238754 75868 240108
rect 74538 238711 74594 238720
rect 74644 238726 75224 238754
rect 75288 238726 75868 238754
rect 73896 238196 73948 238202
rect 73896 238138 73948 238144
rect 73252 237176 73304 237182
rect 73252 237118 73304 237124
rect 73264 236026 73292 237118
rect 73252 236020 73304 236026
rect 73252 235962 73304 235968
rect 73804 236020 73856 236026
rect 73804 235962 73856 235968
rect 73816 185638 73844 235962
rect 74552 204950 74580 238711
rect 74644 215966 74672 238726
rect 75288 233866 75316 238726
rect 75552 237448 75604 237454
rect 75552 237390 75604 237396
rect 74736 233838 75316 233866
rect 74736 229090 74764 233838
rect 75564 233102 75592 237390
rect 76484 233102 76512 240108
rect 77128 237454 77156 240108
rect 77116 237448 77168 237454
rect 77116 237390 77168 237396
rect 75184 233096 75236 233102
rect 75184 233038 75236 233044
rect 75552 233096 75604 233102
rect 75552 233038 75604 233044
rect 76472 233096 76524 233102
rect 76472 233038 76524 233044
rect 74724 229084 74776 229090
rect 74724 229026 74776 229032
rect 74632 215960 74684 215966
rect 74632 215902 74684 215908
rect 74540 204944 74592 204950
rect 74540 204886 74592 204892
rect 73804 185632 73856 185638
rect 73804 185574 73856 185580
rect 75196 184210 75224 233038
rect 77772 233034 77800 240108
rect 78416 238754 78444 240108
rect 78680 238944 78732 238950
rect 78680 238886 78732 238892
rect 77864 238726 78444 238754
rect 77760 233028 77812 233034
rect 77760 232970 77812 232976
rect 77864 219434 77892 238726
rect 77944 233028 77996 233034
rect 77944 232970 77996 232976
rect 77312 219406 77892 219434
rect 77312 192642 77340 219406
rect 77956 198014 77984 232970
rect 78692 211886 78720 238886
rect 79060 222902 79088 240108
rect 79704 238950 79732 240108
rect 79692 238944 79744 238950
rect 79692 238886 79744 238892
rect 80348 235822 80376 240108
rect 80992 238754 81020 240108
rect 81440 239080 81492 239086
rect 81440 239022 81492 239028
rect 80624 238726 81020 238754
rect 80336 235816 80388 235822
rect 80336 235758 80388 235764
rect 80348 234666 80376 235758
rect 80336 234660 80388 234666
rect 80336 234602 80388 234608
rect 79048 222896 79100 222902
rect 79048 222838 79100 222844
rect 80624 219434 80652 238726
rect 80704 234660 80756 234666
rect 80704 234602 80756 234608
rect 80072 219406 80652 219434
rect 78680 211880 78732 211886
rect 78680 211822 78732 211828
rect 80072 208282 80100 219406
rect 80060 208276 80112 208282
rect 80060 208218 80112 208224
rect 77944 198008 77996 198014
rect 77944 197950 77996 197956
rect 77300 192636 77352 192642
rect 77300 192578 77352 192584
rect 80716 185609 80744 234602
rect 81452 224942 81480 239022
rect 81636 237250 81664 240108
rect 82280 239086 82308 240108
rect 82924 239154 82952 240108
rect 82912 239148 82964 239154
rect 82912 239090 82964 239096
rect 82268 239080 82320 239086
rect 82268 239022 82320 239028
rect 82924 238746 82952 239090
rect 83568 238754 83596 240108
rect 82912 238740 82964 238746
rect 82912 238682 82964 238688
rect 83476 238726 83596 238754
rect 84212 238754 84240 240108
rect 84212 238726 84332 238754
rect 81624 237244 81676 237250
rect 81624 237186 81676 237192
rect 81636 231742 81664 237186
rect 83476 234394 83504 238726
rect 83464 234388 83516 234394
rect 83464 234330 83516 234336
rect 81624 231736 81676 231742
rect 81624 231678 81676 231684
rect 81440 224936 81492 224942
rect 81440 224878 81492 224884
rect 83476 213246 83504 234330
rect 84200 233912 84252 233918
rect 84200 233854 84252 233860
rect 83464 213240 83516 213246
rect 83464 213182 83516 213188
rect 84212 209710 84240 233854
rect 84304 213926 84332 238726
rect 84856 233918 84884 240108
rect 84844 233912 84896 233918
rect 84844 233854 84896 233860
rect 85500 222873 85528 240108
rect 86144 238649 86172 240108
rect 86788 238754 86816 240108
rect 86788 238726 86908 238754
rect 86130 238640 86186 238649
rect 86130 238575 86186 238584
rect 86224 238128 86276 238134
rect 86224 238070 86276 238076
rect 85486 222864 85542 222873
rect 85486 222799 85542 222808
rect 84292 213920 84344 213926
rect 84292 213862 84344 213868
rect 84200 209704 84252 209710
rect 84200 209646 84252 209652
rect 86236 209098 86264 238070
rect 86880 234462 86908 238726
rect 87432 235414 87460 240108
rect 88076 238406 88104 240108
rect 88064 238400 88116 238406
rect 88064 238342 88116 238348
rect 88248 235816 88300 235822
rect 88248 235758 88300 235764
rect 88260 235414 88288 235758
rect 87420 235408 87472 235414
rect 87420 235350 87472 235356
rect 88248 235408 88300 235414
rect 88248 235350 88300 235356
rect 86868 234456 86920 234462
rect 86868 234398 86920 234404
rect 86880 233034 86908 234398
rect 86868 233028 86920 233034
rect 86868 232970 86920 232976
rect 86224 209092 86276 209098
rect 86224 209034 86276 209040
rect 88260 189786 88288 235350
rect 88720 231538 88748 240108
rect 89364 238678 89392 240108
rect 89352 238672 89404 238678
rect 89352 238614 89404 238620
rect 89720 233912 89772 233918
rect 89720 233854 89772 233860
rect 88708 231532 88760 231538
rect 88708 231474 88760 231480
rect 89732 210594 89760 233854
rect 90008 220182 90036 240108
rect 90652 233918 90680 240108
rect 91296 238610 91324 240108
rect 91940 238678 91968 240108
rect 91928 238672 91980 238678
rect 91928 238614 91980 238620
rect 91284 238604 91336 238610
rect 91284 238546 91336 238552
rect 91744 238400 91796 238406
rect 91744 238342 91796 238348
rect 90640 233912 90692 233918
rect 90640 233854 90692 233860
rect 89996 220176 90048 220182
rect 89996 220118 90048 220124
rect 89720 210588 89772 210594
rect 89720 210530 89772 210536
rect 91756 195430 91784 238342
rect 92480 238060 92532 238066
rect 92480 238002 92532 238008
rect 92492 237522 92520 238002
rect 92480 237516 92532 237522
rect 92480 237458 92532 237464
rect 92584 219434 92612 240108
rect 93228 238134 93256 240108
rect 93872 238754 93900 240108
rect 93872 238726 94084 238754
rect 93216 238128 93268 238134
rect 93216 238070 93268 238076
rect 93768 237516 93820 237522
rect 93768 237458 93820 237464
rect 92492 219406 92612 219434
rect 92492 203658 92520 219406
rect 92480 203652 92532 203658
rect 92480 203594 92532 203600
rect 93780 199442 93808 237458
rect 93952 233912 94004 233918
rect 93952 233854 94004 233860
rect 93964 216578 93992 233854
rect 93952 216572 94004 216578
rect 93952 216514 94004 216520
rect 93768 199436 93820 199442
rect 93768 199378 93820 199384
rect 91744 195424 91796 195430
rect 91744 195366 91796 195372
rect 88248 189780 88300 189786
rect 88248 189722 88300 189728
rect 80702 185600 80758 185609
rect 80702 185535 80758 185544
rect 75184 184204 75236 184210
rect 75184 184146 75236 184152
rect 73068 182844 73120 182850
rect 73068 182786 73120 182792
rect 94056 181626 94084 238726
rect 94516 233918 94544 240108
rect 95160 237522 95188 240108
rect 95148 237516 95200 237522
rect 95148 237458 95200 237464
rect 95804 237250 95832 240108
rect 96448 239442 96476 240108
rect 96448 239414 96568 239442
rect 96436 239284 96488 239290
rect 96436 239226 96488 239232
rect 95792 237244 95844 237250
rect 95792 237186 95844 237192
rect 94504 233912 94556 233918
rect 94504 233854 94556 233860
rect 96448 205630 96476 239226
rect 96540 238338 96568 239414
rect 96528 238332 96580 238338
rect 96528 238274 96580 238280
rect 96436 205624 96488 205630
rect 96436 205566 96488 205572
rect 96540 186998 96568 238274
rect 97092 219434 97120 240108
rect 97736 239290 97764 240108
rect 97724 239284 97776 239290
rect 97724 239226 97776 239232
rect 98380 230382 98408 240108
rect 99024 238542 99052 240108
rect 99668 238950 99696 240108
rect 99380 238944 99432 238950
rect 99380 238886 99432 238892
rect 99656 238944 99708 238950
rect 99656 238886 99708 238892
rect 99012 238536 99064 238542
rect 99012 238478 99064 238484
rect 98828 238128 98880 238134
rect 98828 238070 98880 238076
rect 98840 237182 98868 238070
rect 98828 237176 98880 237182
rect 98828 237118 98880 237124
rect 99288 237176 99340 237182
rect 99288 237118 99340 237124
rect 98368 230376 98420 230382
rect 98368 230318 98420 230324
rect 96632 219406 97120 219434
rect 96632 196790 96660 219406
rect 96620 196784 96672 196790
rect 96620 196726 96672 196732
rect 99300 194070 99328 237118
rect 99392 202162 99420 238886
rect 100312 219434 100340 240108
rect 100760 233912 100812 233918
rect 100760 233854 100812 233860
rect 99484 219406 100340 219434
rect 99484 218890 99512 219406
rect 99472 218884 99524 218890
rect 99472 218826 99524 218832
rect 99380 202156 99432 202162
rect 99380 202098 99432 202104
rect 99288 194064 99340 194070
rect 99288 194006 99340 194012
rect 100772 192710 100800 233854
rect 100956 227186 100984 240108
rect 101600 233918 101628 240108
rect 102244 235346 102272 240108
rect 102232 235340 102284 235346
rect 102232 235282 102284 235288
rect 101588 233912 101640 233918
rect 101588 233854 101640 233860
rect 100944 227180 100996 227186
rect 100944 227122 100996 227128
rect 102888 219434 102916 240108
rect 103532 237454 103560 240108
rect 103520 237448 103572 237454
rect 103520 237390 103572 237396
rect 103704 233912 103756 233918
rect 103704 233854 103756 233860
rect 102152 219406 102916 219434
rect 100760 192704 100812 192710
rect 100760 192646 100812 192652
rect 102152 189922 102180 219406
rect 103716 215286 103744 233854
rect 104176 230450 104204 240108
rect 104532 237448 104584 237454
rect 104532 237390 104584 237396
rect 104624 237448 104676 237454
rect 104624 237390 104676 237396
rect 104256 231668 104308 231674
rect 104256 231610 104308 231616
rect 104164 230444 104216 230450
rect 104164 230386 104216 230392
rect 103704 215280 103756 215286
rect 103704 215222 103756 215228
rect 104176 192574 104204 230386
rect 104268 206310 104296 231610
rect 104544 230450 104572 237390
rect 104636 231674 104664 237390
rect 104820 233918 104848 240108
rect 105464 238610 105492 240108
rect 105452 238604 105504 238610
rect 105452 238546 105504 238552
rect 106108 237454 106136 240108
rect 106096 237448 106148 237454
rect 106096 237390 106148 237396
rect 106752 237318 106780 240108
rect 107396 239018 107424 240108
rect 107384 239012 107436 239018
rect 107384 238954 107436 238960
rect 108040 237998 108068 240108
rect 108028 237992 108080 237998
rect 108028 237934 108080 237940
rect 106740 237312 106792 237318
rect 106740 237254 106792 237260
rect 104808 233912 104860 233918
rect 104808 233854 104860 233860
rect 104624 231668 104676 231674
rect 104624 231610 104676 231616
rect 104532 230444 104584 230450
rect 104532 230386 104584 230392
rect 108684 227662 108712 240108
rect 109972 238785 110000 240108
rect 109038 238776 109094 238785
rect 109038 238711 109094 238720
rect 109958 238776 110014 238785
rect 109958 238711 110014 238720
rect 108948 238400 109000 238406
rect 108948 238342 109000 238348
rect 108960 237998 108988 238342
rect 108948 237992 109000 237998
rect 108948 237934 109000 237940
rect 108672 227656 108724 227662
rect 108672 227598 108724 227604
rect 108960 214606 108988 237934
rect 108948 214600 109000 214606
rect 108948 214542 109000 214548
rect 104256 206304 104308 206310
rect 104256 206246 104308 206252
rect 104164 192568 104216 192574
rect 104164 192510 104216 192516
rect 102140 189916 102192 189922
rect 102140 189858 102192 189864
rect 109052 189854 109080 238711
rect 110616 234462 110644 240108
rect 111260 239442 111288 240108
rect 110984 239414 111288 239442
rect 110604 234456 110656 234462
rect 110604 234398 110656 234404
rect 110984 219434 111012 239414
rect 111154 239320 111210 239329
rect 111154 239255 111210 239264
rect 111064 234456 111116 234462
rect 111064 234398 111116 234404
rect 110432 219406 111012 219434
rect 110432 203726 110460 219406
rect 110420 203720 110472 203726
rect 110420 203662 110472 203668
rect 109040 189848 109092 189854
rect 109040 189790 109092 189796
rect 106188 189168 106240 189174
rect 106188 189110 106240 189116
rect 102048 187740 102100 187746
rect 102048 187682 102100 187688
rect 96528 186992 96580 186998
rect 96528 186934 96580 186940
rect 100668 185020 100720 185026
rect 100668 184962 100720 184968
rect 94044 181620 94096 181626
rect 94044 181562 94096 181568
rect 68926 181384 68982 181393
rect 68926 181319 68982 181328
rect 64788 180124 64840 180130
rect 64788 180066 64840 180072
rect 100680 177585 100708 184962
rect 102060 177585 102088 187682
rect 104808 186380 104860 186386
rect 104808 186322 104860 186328
rect 104820 177585 104848 186322
rect 106200 177585 106228 189110
rect 109960 177948 110012 177954
rect 109960 177890 110012 177896
rect 100666 177576 100722 177585
rect 100666 177511 100722 177520
rect 102046 177576 102102 177585
rect 102046 177511 102102 177520
rect 104806 177576 104862 177585
rect 104806 177511 104862 177520
rect 106186 177576 106242 177585
rect 106186 177511 106242 177520
rect 108120 176860 108172 176866
rect 108120 176802 108172 176808
rect 107016 176792 107068 176798
rect 107014 176760 107016 176769
rect 108132 176769 108160 176802
rect 109972 176769 110000 177890
rect 107068 176760 107070 176769
rect 107014 176695 107070 176704
rect 108118 176760 108174 176769
rect 108118 176695 108174 176704
rect 109958 176760 110014 176769
rect 109958 176695 110014 176704
rect 98368 176112 98420 176118
rect 98368 176054 98420 176060
rect 98380 175409 98408 176054
rect 100760 176044 100812 176050
rect 100760 175986 100812 175992
rect 100772 175409 100800 175986
rect 111076 175982 111104 234398
rect 111168 184346 111196 239255
rect 111904 219434 111932 240108
rect 112548 235890 112576 240108
rect 112536 235884 112588 235890
rect 112536 235826 112588 235832
rect 113192 232966 113220 240108
rect 113836 233170 113864 240108
rect 114480 237017 114508 240108
rect 114466 237008 114522 237017
rect 114466 236943 114522 236952
rect 114560 233912 114612 233918
rect 114560 233854 114612 233860
rect 114468 233300 114520 233306
rect 114468 233242 114520 233248
rect 113824 233164 113876 233170
rect 113824 233106 113876 233112
rect 114480 232966 114508 233242
rect 113180 232960 113232 232966
rect 113180 232902 113232 232908
rect 114468 232960 114520 232966
rect 114468 232902 114520 232908
rect 111812 219406 111932 219434
rect 111812 213314 111840 219406
rect 111800 213308 111852 213314
rect 111800 213250 111852 213256
rect 114572 208350 114600 233854
rect 115124 231606 115152 240108
rect 115768 233918 115796 240108
rect 115756 233912 115808 233918
rect 115756 233854 115808 233860
rect 115112 231600 115164 231606
rect 115112 231542 115164 231548
rect 116412 219434 116440 240108
rect 117056 239902 117084 240108
rect 117044 239896 117096 239902
rect 117044 239838 117096 239844
rect 117700 238513 117728 240108
rect 117686 238504 117742 238513
rect 117686 238439 117688 238448
rect 117740 238439 117742 238448
rect 117688 238410 117740 238416
rect 117700 238379 117728 238410
rect 117964 233300 118016 233306
rect 117964 233242 118016 233248
rect 115952 219406 116440 219434
rect 114560 208344 114612 208350
rect 114560 208286 114612 208292
rect 115952 207806 115980 219406
rect 115940 207800 115992 207806
rect 115940 207742 115992 207748
rect 117976 195265 118004 233242
rect 118344 230314 118372 240108
rect 118988 239970 119016 240108
rect 119646 240094 119844 240122
rect 118976 239964 119028 239970
rect 118976 239906 119028 239912
rect 119816 238746 119844 240094
rect 119908 239970 119936 240887
rect 119896 239964 119948 239970
rect 119896 239906 119948 239912
rect 120000 238754 120028 242218
rect 120078 241496 120134 241505
rect 120078 241431 120134 241440
rect 119804 238740 119856 238746
rect 119804 238682 119856 238688
rect 119908 238726 120028 238754
rect 118332 230308 118384 230314
rect 118332 230250 118384 230256
rect 119816 229094 119844 238682
rect 119908 238338 119936 238726
rect 119896 238332 119948 238338
rect 119896 238274 119948 238280
rect 119816 229066 120028 229094
rect 120000 202298 120028 229066
rect 119988 202292 120040 202298
rect 119988 202234 120040 202240
rect 117962 195256 118018 195265
rect 117962 195191 118018 195200
rect 111156 184340 111208 184346
rect 111156 184282 111208 184288
rect 118424 182232 118476 182238
rect 114006 182200 114062 182209
rect 118424 182174 118476 182180
rect 114006 182135 114062 182144
rect 112444 178288 112496 178294
rect 112444 178230 112496 178236
rect 112456 176769 112484 178230
rect 114020 177585 114048 182135
rect 114284 179444 114336 179450
rect 114284 179386 114336 179392
rect 114006 177576 114062 177585
rect 114006 177511 114062 177520
rect 114296 177041 114324 179386
rect 118436 177585 118464 182174
rect 120092 178022 120120 241431
rect 120184 224262 120212 250951
rect 120736 239902 120764 253914
rect 120828 244934 120856 291858
rect 121472 291825 121500 383658
rect 121552 309800 121604 309806
rect 121552 309742 121604 309748
rect 121458 291816 121514 291825
rect 121458 291751 121514 291760
rect 121458 290456 121514 290465
rect 121458 290391 121514 290400
rect 121472 290018 121500 290391
rect 121460 290012 121512 290018
rect 121460 289954 121512 289960
rect 121460 289808 121512 289814
rect 121460 289750 121512 289756
rect 121472 289105 121500 289750
rect 121458 289096 121514 289105
rect 121458 289031 121514 289040
rect 121460 288380 121512 288386
rect 121460 288322 121512 288328
rect 121472 287745 121500 288322
rect 121458 287736 121514 287745
rect 121458 287671 121514 287680
rect 121564 285818 121592 309742
rect 122116 306374 122144 402222
rect 123956 401674 123984 405076
rect 124220 403640 124272 403646
rect 124220 403582 124272 403588
rect 123944 401668 123996 401674
rect 123944 401610 123996 401616
rect 123484 398200 123536 398206
rect 123484 398142 123536 398148
rect 122748 360868 122800 360874
rect 122748 360810 122800 360816
rect 122116 306346 122236 306374
rect 121642 291136 121698 291145
rect 121642 291071 121698 291080
rect 121656 289950 121684 291071
rect 121644 289944 121696 289950
rect 121644 289886 121696 289892
rect 121642 288416 121698 288425
rect 121642 288351 121698 288360
rect 121656 287094 121684 288351
rect 121644 287088 121696 287094
rect 121644 287030 121696 287036
rect 121564 285790 121684 285818
rect 121552 285660 121604 285666
rect 121552 285602 121604 285608
rect 121460 285592 121512 285598
rect 121460 285534 121512 285540
rect 121472 285025 121500 285534
rect 121458 285016 121514 285025
rect 121458 284951 121514 284960
rect 121564 284345 121592 285602
rect 121550 284336 121606 284345
rect 121550 284271 121606 284280
rect 121458 282976 121514 282985
rect 121458 282911 121460 282920
rect 121512 282911 121514 282920
rect 121460 282882 121512 282888
rect 121550 282296 121606 282305
rect 121550 282231 121606 282240
rect 121564 281654 121592 282231
rect 121552 281648 121604 281654
rect 121458 281616 121514 281625
rect 121552 281590 121604 281596
rect 121458 281551 121460 281560
rect 121512 281551 121514 281560
rect 121460 281522 121512 281528
rect 121458 280256 121514 280265
rect 121458 280191 121460 280200
rect 121512 280191 121514 280200
rect 121460 280162 121512 280168
rect 121458 278896 121514 278905
rect 121458 278831 121514 278840
rect 121472 278798 121500 278831
rect 121460 278792 121512 278798
rect 121656 278769 121684 285790
rect 122208 284986 122236 306346
rect 122196 284980 122248 284986
rect 122196 284922 122248 284928
rect 122102 280936 122158 280945
rect 122102 280871 122158 280880
rect 121460 278734 121512 278740
rect 121642 278760 121698 278769
rect 121552 278724 121604 278730
rect 121642 278695 121698 278704
rect 121552 278666 121604 278672
rect 121564 277545 121592 278666
rect 121550 277536 121606 277545
rect 121550 277471 121606 277480
rect 121460 277364 121512 277370
rect 121460 277306 121512 277312
rect 121472 276865 121500 277306
rect 121458 276856 121514 276865
rect 121458 276791 121514 276800
rect 121458 275496 121514 275505
rect 121458 275431 121514 275440
rect 121472 274786 121500 275431
rect 121550 274816 121606 274825
rect 121460 274780 121512 274786
rect 121550 274751 121606 274760
rect 121460 274722 121512 274728
rect 121564 274718 121592 274751
rect 121552 274712 121604 274718
rect 121552 274654 121604 274660
rect 121460 274644 121512 274650
rect 121460 274586 121512 274592
rect 121472 274145 121500 274586
rect 121458 274136 121514 274145
rect 121458 274071 121514 274080
rect 121458 273456 121514 273465
rect 121458 273391 121514 273400
rect 121472 273290 121500 273391
rect 121460 273284 121512 273290
rect 121460 273226 121512 273232
rect 121458 272776 121514 272785
rect 121458 272711 121514 272720
rect 121472 272610 121500 272711
rect 121460 272604 121512 272610
rect 121460 272546 121512 272552
rect 121458 271416 121514 271425
rect 121458 271351 121514 271360
rect 121472 270570 121500 271351
rect 121460 270564 121512 270570
rect 121460 270506 121512 270512
rect 121458 270056 121514 270065
rect 121458 269991 121514 270000
rect 120908 269816 120960 269822
rect 120908 269758 120960 269764
rect 120816 244928 120868 244934
rect 120816 244870 120868 244876
rect 120724 239896 120776 239902
rect 120724 239838 120776 239844
rect 120920 238542 120948 269758
rect 121472 269210 121500 269991
rect 121550 269376 121606 269385
rect 121550 269311 121606 269320
rect 121460 269204 121512 269210
rect 121460 269146 121512 269152
rect 121564 269142 121592 269311
rect 121552 269136 121604 269142
rect 121552 269078 121604 269084
rect 121460 269068 121512 269074
rect 121460 269010 121512 269016
rect 121472 268705 121500 269010
rect 121458 268696 121514 268705
rect 121458 268631 121514 268640
rect 121460 268388 121512 268394
rect 121460 268330 121512 268336
rect 121472 268025 121500 268330
rect 121458 268016 121514 268025
rect 121458 267951 121514 267960
rect 121552 267708 121604 267714
rect 121552 267650 121604 267656
rect 121458 267336 121514 267345
rect 121458 267271 121514 267280
rect 121472 266422 121500 267271
rect 121564 266665 121592 267650
rect 121550 266656 121606 266665
rect 121550 266591 121606 266600
rect 121460 266416 121512 266422
rect 121460 266358 121512 266364
rect 121458 264616 121514 264625
rect 121458 264551 121514 264560
rect 121472 264246 121500 264551
rect 121460 264240 121512 264246
rect 121460 264182 121512 264188
rect 121550 263936 121606 263945
rect 121550 263871 121606 263880
rect 121564 263634 121592 263871
rect 121552 263628 121604 263634
rect 121552 263570 121604 263576
rect 121460 263560 121512 263566
rect 121460 263502 121512 263508
rect 121472 263265 121500 263502
rect 121458 263256 121514 263265
rect 121458 263191 121514 263200
rect 121460 262880 121512 262886
rect 121460 262822 121512 262828
rect 121472 262585 121500 262822
rect 121458 262576 121514 262585
rect 121458 262511 121514 262520
rect 121000 262268 121052 262274
rect 121000 262210 121052 262216
rect 121012 261905 121040 262210
rect 121460 262200 121512 262206
rect 121460 262142 121512 262148
rect 120998 261896 121054 261905
rect 120998 261831 121054 261840
rect 121472 261225 121500 262142
rect 121458 261216 121514 261225
rect 121458 261151 121514 261160
rect 121460 260840 121512 260846
rect 121460 260782 121512 260788
rect 121472 260545 121500 260782
rect 121458 260536 121514 260545
rect 121458 260471 121514 260480
rect 122116 260166 122144 280871
rect 122760 279585 122788 360810
rect 122840 284980 122892 284986
rect 122840 284922 122892 284928
rect 122746 279576 122802 279585
rect 122746 279511 122802 279520
rect 122760 279478 122788 279511
rect 122748 279472 122800 279478
rect 122748 279414 122800 279420
rect 122286 278760 122342 278769
rect 122286 278695 122342 278704
rect 122194 265976 122250 265985
rect 122194 265911 122250 265920
rect 122104 260160 122156 260166
rect 122104 260102 122156 260108
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259486 121500 259791
rect 121460 259480 121512 259486
rect 121460 259422 121512 259428
rect 122102 259176 122158 259185
rect 122102 259111 122158 259120
rect 121458 258496 121514 258505
rect 121458 258431 121514 258440
rect 121472 258126 121500 258431
rect 121460 258120 121512 258126
rect 121460 258062 121512 258068
rect 121550 257816 121606 257825
rect 121550 257751 121606 257760
rect 121458 257136 121514 257145
rect 121458 257071 121514 257080
rect 121472 256834 121500 257071
rect 121564 256902 121592 257751
rect 121552 256896 121604 256902
rect 121552 256838 121604 256844
rect 121460 256828 121512 256834
rect 121460 256770 121512 256776
rect 121550 256456 121606 256465
rect 121550 256391 121606 256400
rect 121458 255776 121514 255785
rect 121458 255711 121514 255720
rect 121472 255338 121500 255711
rect 121564 255406 121592 256391
rect 121552 255400 121604 255406
rect 121552 255342 121604 255348
rect 121460 255332 121512 255338
rect 121460 255274 121512 255280
rect 121458 254416 121514 254425
rect 121458 254351 121514 254360
rect 121472 254046 121500 254351
rect 121460 254040 121512 254046
rect 121460 253982 121512 253988
rect 121460 253904 121512 253910
rect 121460 253846 121512 253852
rect 121472 253065 121500 253846
rect 121550 253736 121606 253745
rect 121550 253671 121606 253680
rect 121458 253056 121514 253065
rect 121458 252991 121514 253000
rect 121564 252618 121592 253671
rect 121552 252612 121604 252618
rect 121552 252554 121604 252560
rect 121458 252376 121514 252385
rect 121458 252311 121514 252320
rect 121472 251258 121500 252311
rect 121460 251252 121512 251258
rect 121460 251194 121512 251200
rect 121550 250336 121606 250345
rect 121550 250271 121606 250280
rect 121564 249830 121592 250271
rect 121552 249824 121604 249830
rect 121552 249766 121604 249772
rect 121460 249756 121512 249762
rect 121460 249698 121512 249704
rect 121472 249665 121500 249698
rect 121458 249656 121514 249665
rect 121458 249591 121514 249600
rect 121460 248396 121512 248402
rect 121460 248338 121512 248344
rect 121472 247625 121500 248338
rect 121550 248296 121606 248305
rect 121550 248231 121606 248240
rect 121458 247616 121514 247625
rect 121458 247551 121514 247560
rect 121564 247110 121592 248231
rect 121552 247104 121604 247110
rect 121552 247046 121604 247052
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 121458 246256 121514 246265
rect 121458 246191 121514 246200
rect 121472 245682 121500 246191
rect 121564 245750 121592 246871
rect 121552 245744 121604 245750
rect 121552 245686 121604 245692
rect 121460 245676 121512 245682
rect 121460 245618 121512 245624
rect 121552 245608 121604 245614
rect 121458 245576 121514 245585
rect 121552 245550 121604 245556
rect 121458 245511 121514 245520
rect 121472 245070 121500 245511
rect 121460 245064 121512 245070
rect 121460 245006 121512 245012
rect 121564 244905 121592 245550
rect 121550 244896 121606 244905
rect 121550 244831 121606 244840
rect 121460 244248 121512 244254
rect 121458 244216 121460 244225
rect 121512 244216 121514 244225
rect 121458 244151 121514 244160
rect 121552 242888 121604 242894
rect 121458 242856 121514 242865
rect 121552 242830 121604 242836
rect 121458 242791 121460 242800
rect 121512 242791 121514 242800
rect 121460 242762 121512 242768
rect 121564 242185 121592 242830
rect 121550 242176 121606 242185
rect 121550 242111 121606 242120
rect 121458 240816 121514 240825
rect 121458 240751 121514 240760
rect 121472 240174 121500 240751
rect 121460 240168 121512 240174
rect 121460 240110 121512 240116
rect 121550 240136 121606 240145
rect 121550 240071 121606 240080
rect 121564 240038 121592 240071
rect 121552 240032 121604 240038
rect 121552 239974 121604 239980
rect 120908 238536 120960 238542
rect 120908 238478 120960 238484
rect 122116 228993 122144 259111
rect 122208 258074 122236 265911
rect 122300 258738 122328 278695
rect 122378 272096 122434 272105
rect 122378 272031 122434 272040
rect 122392 267734 122420 272031
rect 122392 267706 122512 267734
rect 122288 258732 122340 258738
rect 122288 258674 122340 258680
rect 122208 258046 122328 258074
rect 122194 251696 122250 251705
rect 122194 251631 122250 251640
rect 122102 228984 122158 228993
rect 122102 228919 122158 228928
rect 120172 224256 120224 224262
rect 120172 224198 120224 224204
rect 122104 220244 122156 220250
rect 122104 220186 122156 220192
rect 122116 182918 122144 220186
rect 122208 216646 122236 251631
rect 122300 238066 122328 258046
rect 122484 256018 122512 267706
rect 122472 256012 122524 256018
rect 122472 255954 122524 255960
rect 122378 255096 122434 255105
rect 122378 255031 122434 255040
rect 122392 248414 122420 255031
rect 122392 248386 122512 248414
rect 122288 238060 122340 238066
rect 122288 238002 122340 238008
rect 122484 237386 122512 248386
rect 122472 237380 122524 237386
rect 122472 237322 122524 237328
rect 122196 216640 122248 216646
rect 122196 216582 122248 216588
rect 122852 208282 122880 284922
rect 122930 248976 122986 248985
rect 122930 248911 122986 248920
rect 122944 229022 122972 248911
rect 123496 238406 123524 398142
rect 123668 294228 123720 294234
rect 123668 294170 123720 294176
rect 123680 280838 123708 294170
rect 123760 292868 123812 292874
rect 123760 292810 123812 292816
rect 123772 282878 123800 292810
rect 123760 282872 123812 282878
rect 123760 282814 123812 282820
rect 123668 280832 123720 280838
rect 123668 280774 123720 280780
rect 124232 272610 124260 403582
rect 126980 402348 127032 402354
rect 126980 402290 127032 402296
rect 124864 393984 124916 393990
rect 124864 393926 124916 393932
rect 124312 311228 124364 311234
rect 124312 311170 124364 311176
rect 124220 272604 124272 272610
rect 124220 272546 124272 272552
rect 124324 262886 124352 311170
rect 124402 286648 124458 286657
rect 124402 286583 124458 286592
rect 124416 285734 124444 286583
rect 124404 285728 124456 285734
rect 124404 285670 124456 285676
rect 124312 262880 124364 262886
rect 124312 262822 124364 262828
rect 123576 256760 123628 256766
rect 123576 256702 123628 256708
rect 123484 238400 123536 238406
rect 123484 238342 123536 238348
rect 123588 237318 123616 256702
rect 124876 238746 124904 393926
rect 126244 381540 126296 381546
rect 126244 381482 126296 381488
rect 124956 294160 125008 294166
rect 124956 294102 125008 294108
rect 124864 238740 124916 238746
rect 124864 238682 124916 238688
rect 123576 237312 123628 237318
rect 123576 237254 123628 237260
rect 122932 229016 122984 229022
rect 122932 228958 122984 228964
rect 122944 227798 122972 228958
rect 122932 227792 122984 227798
rect 122932 227734 122984 227740
rect 124864 227792 124916 227798
rect 124864 227734 124916 227740
rect 122840 208276 122892 208282
rect 122840 208218 122892 208224
rect 124128 208276 124180 208282
rect 124128 208218 124180 208224
rect 124140 207738 124168 208218
rect 124128 207732 124180 207738
rect 124128 207674 124180 207680
rect 124876 191418 124904 227734
rect 124968 194002 124996 294102
rect 126256 268394 126284 381482
rect 126888 341556 126940 341562
rect 126888 341498 126940 341504
rect 126900 341465 126928 341498
rect 126886 341456 126942 341465
rect 126886 341391 126942 341400
rect 126428 314016 126480 314022
rect 126428 313958 126480 313964
rect 126336 295588 126388 295594
rect 126336 295530 126388 295536
rect 126244 268388 126296 268394
rect 126244 268330 126296 268336
rect 126256 198082 126284 268330
rect 126348 209234 126376 295530
rect 126440 289814 126468 313958
rect 126520 292936 126572 292942
rect 126520 292878 126572 292884
rect 126428 289808 126480 289814
rect 126428 289750 126480 289756
rect 126428 287700 126480 287706
rect 126428 287642 126480 287648
rect 126440 237182 126468 287642
rect 126532 276010 126560 292878
rect 126520 276004 126572 276010
rect 126520 275946 126572 275952
rect 126428 237176 126480 237182
rect 126428 237118 126480 237124
rect 126992 235822 127020 402290
rect 127176 401674 127204 405076
rect 129752 405062 130410 405090
rect 132512 405062 133630 405090
rect 127164 401668 127216 401674
rect 127164 401610 127216 401616
rect 129004 401668 129056 401674
rect 129004 401610 129056 401616
rect 127808 308440 127860 308446
rect 127808 308382 127860 308388
rect 127624 295656 127676 295662
rect 127624 295598 127676 295604
rect 127532 238740 127584 238746
rect 127532 238682 127584 238688
rect 127544 238474 127572 238682
rect 127532 238468 127584 238474
rect 127532 238410 127584 238416
rect 126980 235816 127032 235822
rect 126980 235758 127032 235764
rect 126336 209228 126388 209234
rect 126336 209170 126388 209176
rect 126244 198076 126296 198082
rect 126244 198018 126296 198024
rect 124956 193996 125008 194002
rect 124956 193938 125008 193944
rect 124864 191412 124916 191418
rect 124864 191354 124916 191360
rect 127636 188426 127664 295598
rect 127716 291848 127768 291854
rect 127716 291790 127768 291796
rect 127728 242826 127756 291790
rect 127820 277370 127848 308382
rect 127808 277364 127860 277370
rect 127808 277306 127860 277312
rect 128360 272536 128412 272542
rect 128360 272478 128412 272484
rect 128372 269822 128400 272478
rect 128360 269816 128412 269822
rect 128360 269758 128412 269764
rect 128360 247036 128412 247042
rect 128360 246978 128412 246984
rect 127716 242820 127768 242826
rect 127716 242762 127768 242768
rect 128372 240961 128400 246978
rect 128358 240952 128414 240961
rect 128358 240887 128414 240896
rect 129016 231878 129044 401610
rect 129752 367810 129780 405062
rect 132408 384328 132460 384334
rect 132408 384270 132460 384276
rect 129832 371884 129884 371890
rect 129832 371826 129884 371832
rect 129844 371278 129872 371826
rect 129832 371272 129884 371278
rect 129832 371214 129884 371220
rect 129740 367804 129792 367810
rect 129740 367746 129792 367752
rect 129096 358896 129148 358902
rect 129096 358838 129148 358844
rect 129108 234462 129136 358838
rect 129280 297424 129332 297430
rect 129280 297366 129332 297372
rect 129188 291236 129240 291242
rect 129188 291178 129240 291184
rect 129096 234456 129148 234462
rect 129096 234398 129148 234404
rect 128360 231872 128412 231878
rect 128360 231814 128412 231820
rect 129004 231872 129056 231878
rect 129004 231814 129056 231820
rect 128372 231538 128400 231814
rect 128360 231532 128412 231538
rect 128360 231474 128412 231480
rect 129200 204921 129228 291178
rect 129292 272542 129320 297366
rect 129740 278724 129792 278730
rect 129740 278666 129792 278672
rect 129752 278050 129780 278666
rect 129740 278044 129792 278050
rect 129740 277986 129792 277992
rect 129280 272536 129332 272542
rect 129280 272478 129332 272484
rect 129844 263566 129872 371214
rect 131026 362264 131082 362273
rect 131026 362199 131082 362208
rect 130476 319456 130528 319462
rect 130476 319398 130528 319404
rect 129832 263560 129884 263566
rect 129832 263502 129884 263508
rect 130384 256012 130436 256018
rect 130384 255954 130436 255960
rect 129648 235408 129700 235414
rect 129648 235350 129700 235356
rect 129660 210526 129688 235350
rect 129648 210520 129700 210526
rect 129648 210462 129700 210468
rect 129186 204912 129242 204921
rect 129186 204847 129242 204856
rect 127624 188420 127676 188426
rect 127624 188362 127676 188368
rect 125508 184952 125560 184958
rect 125508 184894 125560 184900
rect 122104 182912 122156 182918
rect 122104 182854 122156 182860
rect 122012 180872 122064 180878
rect 122012 180814 122064 180820
rect 121000 179580 121052 179586
rect 121000 179522 121052 179528
rect 120080 178016 120132 178022
rect 120080 177958 120132 177964
rect 118422 177576 118478 177585
rect 118422 177511 118478 177520
rect 121012 177041 121040 179522
rect 122024 177585 122052 180814
rect 123024 179648 123076 179654
rect 123024 179590 123076 179596
rect 122010 177576 122066 177585
rect 122010 177511 122066 177520
rect 123036 177041 123064 179590
rect 125520 177585 125548 184894
rect 130396 181665 130424 255954
rect 130488 249762 130516 319398
rect 130568 284980 130620 284986
rect 130568 284922 130620 284928
rect 130476 249756 130528 249762
rect 130476 249698 130528 249704
rect 130580 235414 130608 284922
rect 131040 278050 131068 362199
rect 131120 355360 131172 355366
rect 131120 355302 131172 355308
rect 131132 355094 131160 355302
rect 131120 355088 131172 355094
rect 131120 355030 131172 355036
rect 131028 278044 131080 278050
rect 131028 277986 131080 277992
rect 131132 235890 131160 355030
rect 131856 305108 131908 305114
rect 131856 305050 131908 305056
rect 131764 295520 131816 295526
rect 131764 295462 131816 295468
rect 131212 285796 131264 285802
rect 131212 285738 131264 285744
rect 131224 285598 131252 285738
rect 131212 285592 131264 285598
rect 131212 285534 131264 285540
rect 131120 235884 131172 235890
rect 131120 235826 131172 235832
rect 130568 235408 130620 235414
rect 130568 235350 130620 235356
rect 131776 187202 131804 295462
rect 131868 200870 131896 305050
rect 132420 285802 132448 384270
rect 132512 340950 132540 405062
rect 136836 402286 136864 405076
rect 139412 405062 140070 405090
rect 142172 405062 143290 405090
rect 146312 405062 146510 405090
rect 149072 405062 149730 405090
rect 151832 405062 152950 405090
rect 155972 405062 156170 405090
rect 136824 402280 136876 402286
rect 136824 402222 136876 402228
rect 136640 399560 136692 399566
rect 136640 399502 136692 399508
rect 135904 396976 135956 396982
rect 135904 396918 135956 396924
rect 132590 356144 132646 356153
rect 132590 356079 132646 356088
rect 132500 340944 132552 340950
rect 132500 340886 132552 340892
rect 132500 308508 132552 308514
rect 132500 308450 132552 308456
rect 132408 285796 132460 285802
rect 132408 285738 132460 285744
rect 132512 247042 132540 308450
rect 132604 303006 132632 356079
rect 133972 348424 134024 348430
rect 133972 348366 134024 348372
rect 134616 348424 134668 348430
rect 134616 348366 134668 348372
rect 132868 340944 132920 340950
rect 132868 340886 132920 340892
rect 132880 340202 132908 340886
rect 132868 340196 132920 340202
rect 132868 340138 132920 340144
rect 133880 318164 133932 318170
rect 133880 318106 133932 318112
rect 133144 306468 133196 306474
rect 133144 306410 133196 306416
rect 132592 303000 132644 303006
rect 132592 302942 132644 302948
rect 132500 247036 132552 247042
rect 132500 246978 132552 246984
rect 133156 206378 133184 306410
rect 133236 298376 133288 298382
rect 133236 298318 133288 298324
rect 133144 206372 133196 206378
rect 133144 206314 133196 206320
rect 133248 203794 133276 298318
rect 133892 213926 133920 318106
rect 133984 251190 134012 348366
rect 134628 347818 134656 348366
rect 134616 347812 134668 347818
rect 134616 347754 134668 347760
rect 134524 333260 134576 333266
rect 134524 333202 134576 333208
rect 134536 314090 134564 333202
rect 134524 314084 134576 314090
rect 134524 314026 134576 314032
rect 134616 291304 134668 291310
rect 134616 291246 134668 291252
rect 133972 251184 134024 251190
rect 133972 251126 134024 251132
rect 134524 249824 134576 249830
rect 134524 249766 134576 249772
rect 133880 213920 133932 213926
rect 133880 213862 133932 213868
rect 133236 203788 133288 203794
rect 133236 203730 133288 203736
rect 131856 200864 131908 200870
rect 131856 200806 131908 200812
rect 134536 199578 134564 249766
rect 134628 245002 134656 291246
rect 135168 255400 135220 255406
rect 135168 255342 135220 255348
rect 134616 244996 134668 245002
rect 134616 244938 134668 244944
rect 135180 240786 135208 255342
rect 135168 240780 135220 240786
rect 135168 240722 135220 240728
rect 135916 238950 135944 396918
rect 135996 387932 136048 387938
rect 135996 387874 136048 387880
rect 136008 269074 136036 387874
rect 136088 292732 136140 292738
rect 136088 292674 136140 292680
rect 135996 269068 136048 269074
rect 135996 269010 136048 269016
rect 135904 238944 135956 238950
rect 135904 238886 135956 238892
rect 135168 213920 135220 213926
rect 135168 213862 135220 213868
rect 135180 213246 135208 213862
rect 135168 213240 135220 213246
rect 135168 213182 135220 213188
rect 134524 199572 134576 199578
rect 134524 199514 134576 199520
rect 136100 191350 136128 292674
rect 136180 280220 136232 280226
rect 136180 280162 136232 280168
rect 136192 224262 136220 280162
rect 136180 224256 136232 224262
rect 136180 224198 136232 224204
rect 136652 209710 136680 399502
rect 138020 382968 138072 382974
rect 138020 382910 138072 382916
rect 138032 382294 138060 382910
rect 138020 382288 138072 382294
rect 138020 382230 138072 382236
rect 137284 373312 137336 373318
rect 137284 373254 137336 373260
rect 137296 233102 137324 373254
rect 137376 291372 137428 291378
rect 137376 291314 137428 291320
rect 137284 233096 137336 233102
rect 137284 233038 137336 233044
rect 137388 212022 137416 291314
rect 138032 285666 138060 382230
rect 139308 370524 139360 370530
rect 139308 370466 139360 370472
rect 138664 296812 138716 296818
rect 138664 296754 138716 296760
rect 138020 285660 138072 285666
rect 138020 285602 138072 285608
rect 137376 212016 137428 212022
rect 137376 211958 137428 211964
rect 136640 209704 136692 209710
rect 136640 209646 136692 209652
rect 136652 209166 136680 209646
rect 136640 209160 136692 209166
rect 136640 209102 136692 209108
rect 138676 198150 138704 296754
rect 138756 270564 138808 270570
rect 138756 270506 138808 270512
rect 138664 198144 138716 198150
rect 138664 198086 138716 198092
rect 136088 191344 136140 191350
rect 136088 191286 136140 191292
rect 134524 189100 134576 189106
rect 134524 189042 134576 189048
rect 131764 187196 131816 187202
rect 131764 187138 131816 187144
rect 132408 186448 132460 186454
rect 132408 186390 132460 186396
rect 130382 181656 130438 181665
rect 130382 181591 130438 181600
rect 128176 179512 128228 179518
rect 128176 179454 128228 179460
rect 125506 177576 125562 177585
rect 125506 177511 125562 177520
rect 114282 177032 114338 177041
rect 114282 176967 114338 176976
rect 120998 177032 121054 177041
rect 120998 176967 121054 176976
rect 123022 177032 123078 177041
rect 123022 176967 123078 176976
rect 127072 176996 127124 177002
rect 127072 176938 127124 176944
rect 125784 176928 125836 176934
rect 125784 176870 125836 176876
rect 125796 176769 125824 176870
rect 127084 176769 127112 176938
rect 128188 176769 128216 179454
rect 130752 178220 130804 178226
rect 130752 178162 130804 178168
rect 130764 176769 130792 178162
rect 132420 177585 132448 186390
rect 133604 180940 133656 180946
rect 133604 180882 133656 180888
rect 133616 177585 133644 180882
rect 134536 177954 134564 189042
rect 138768 178702 138796 270506
rect 138848 252612 138900 252618
rect 138848 252554 138900 252560
rect 138860 195498 138888 252554
rect 139320 245818 139348 370466
rect 139412 287706 139440 405062
rect 140780 396772 140832 396778
rect 140780 396714 140832 396720
rect 139490 327720 139546 327729
rect 139490 327655 139546 327664
rect 139504 327146 139532 327655
rect 139492 327140 139544 327146
rect 139492 327082 139544 327088
rect 139400 287700 139452 287706
rect 139400 287642 139452 287648
rect 139308 245812 139360 245818
rect 139308 245754 139360 245760
rect 139504 239018 139532 327082
rect 140136 298172 140188 298178
rect 140136 298114 140188 298120
rect 140044 294024 140096 294030
rect 140044 293966 140096 293972
rect 139492 239012 139544 239018
rect 139492 238954 139544 238960
rect 138848 195492 138900 195498
rect 138848 195434 138900 195440
rect 140056 188494 140084 293966
rect 140148 262138 140176 298114
rect 140228 262880 140280 262886
rect 140228 262822 140280 262828
rect 140136 262132 140188 262138
rect 140136 262074 140188 262080
rect 140136 245812 140188 245818
rect 140136 245754 140188 245760
rect 140148 245070 140176 245754
rect 140136 245064 140188 245070
rect 140136 245006 140188 245012
rect 140148 193866 140176 245006
rect 140240 222970 140268 262822
rect 140792 255406 140820 396714
rect 142172 300830 142200 405062
rect 146312 402974 146340 405062
rect 148416 403640 148468 403646
rect 148416 403582 148468 403588
rect 146220 402946 146340 402974
rect 145564 399492 145616 399498
rect 145564 399434 145616 399440
rect 143540 367804 143592 367810
rect 143540 367746 143592 367752
rect 144276 367804 144328 367810
rect 144276 367746 144328 367752
rect 142896 306400 142948 306406
rect 142896 306342 142948 306348
rect 142160 300824 142212 300830
rect 142160 300766 142212 300772
rect 141514 294128 141570 294137
rect 141514 294063 141570 294072
rect 141424 278792 141476 278798
rect 141424 278734 141476 278740
rect 140780 255400 140832 255406
rect 140780 255342 140832 255348
rect 140228 222964 140280 222970
rect 140228 222906 140280 222912
rect 140136 193860 140188 193866
rect 140136 193802 140188 193808
rect 140044 188488 140096 188494
rect 140044 188430 140096 188436
rect 141436 185774 141464 278734
rect 141528 236706 141556 294063
rect 142802 291952 142858 291961
rect 142802 291887 142858 291896
rect 141608 260160 141660 260166
rect 141608 260102 141660 260108
rect 141516 236700 141568 236706
rect 141516 236642 141568 236648
rect 141620 220250 141648 260102
rect 141608 220244 141660 220250
rect 141608 220186 141660 220192
rect 142816 188465 142844 291887
rect 142908 218822 142936 306342
rect 143448 300824 143500 300830
rect 143448 300766 143500 300772
rect 142988 299804 143040 299810
rect 142988 299746 143040 299752
rect 142896 218816 142948 218822
rect 142896 218758 142948 218764
rect 143000 216170 143028 299746
rect 143460 299538 143488 300766
rect 143448 299532 143500 299538
rect 143448 299474 143500 299480
rect 143460 291854 143488 299474
rect 143448 291848 143500 291854
rect 143448 291790 143500 291796
rect 143552 242894 143580 367746
rect 144288 367130 144316 367746
rect 144276 367124 144328 367130
rect 144276 367066 144328 367072
rect 144184 363656 144236 363662
rect 144184 363598 144236 363604
rect 143632 301572 143684 301578
rect 143632 301514 143684 301520
rect 143644 301481 143672 301514
rect 143630 301472 143686 301481
rect 143630 301407 143686 301416
rect 143540 242888 143592 242894
rect 143540 242830 143592 242836
rect 144196 234394 144224 363598
rect 145576 302326 145604 399434
rect 145564 302320 145616 302326
rect 145564 302262 145616 302268
rect 145748 302320 145800 302326
rect 145748 302262 145800 302268
rect 145564 298240 145616 298246
rect 145564 298182 145616 298188
rect 144276 290012 144328 290018
rect 144276 289954 144328 289960
rect 144184 234388 144236 234394
rect 144184 234330 144236 234336
rect 142988 216164 143040 216170
rect 142988 216106 143040 216112
rect 144288 193934 144316 289954
rect 144368 247104 144420 247110
rect 144368 247046 144420 247052
rect 144380 196926 144408 247046
rect 145576 227254 145604 298182
rect 145656 277432 145708 277438
rect 145656 277374 145708 277380
rect 145668 237318 145696 277374
rect 145760 272649 145788 302262
rect 145746 272640 145802 272649
rect 145746 272575 145802 272584
rect 145656 237312 145708 237318
rect 145656 237254 145708 237260
rect 145564 227248 145616 227254
rect 145564 227190 145616 227196
rect 146220 205630 146248 402946
rect 146300 402280 146352 402286
rect 146300 402222 146352 402228
rect 146312 216578 146340 402222
rect 147586 401024 147642 401033
rect 147586 400959 147642 400968
rect 147128 272604 147180 272610
rect 147128 272546 147180 272552
rect 146944 263628 146996 263634
rect 146944 263570 146996 263576
rect 146300 216572 146352 216578
rect 146300 216514 146352 216520
rect 146312 216034 146340 216514
rect 146300 216028 146352 216034
rect 146300 215970 146352 215976
rect 146208 205624 146260 205630
rect 146208 205566 146260 205572
rect 146220 205086 146248 205566
rect 146208 205080 146260 205086
rect 146208 205022 146260 205028
rect 146956 203862 146984 263570
rect 147036 245744 147088 245750
rect 147036 245686 147088 245692
rect 147048 213382 147076 245686
rect 147140 241233 147168 272546
rect 147600 266257 147628 400959
rect 148324 395344 148376 395350
rect 148324 395286 148376 395292
rect 148336 267714 148364 395286
rect 148428 298314 148456 403582
rect 149072 298761 149100 405062
rect 149704 392012 149756 392018
rect 149704 391954 149756 391960
rect 149058 298752 149114 298761
rect 149058 298687 149114 298696
rect 148416 298308 148468 298314
rect 148416 298250 148468 298256
rect 148324 267708 148376 267714
rect 148324 267650 148376 267656
rect 147586 266248 147642 266257
rect 147586 266183 147642 266192
rect 147600 265577 147628 266183
rect 147586 265568 147642 265577
rect 147586 265503 147642 265512
rect 148324 256896 148376 256902
rect 148324 256838 148376 256844
rect 147126 241224 147182 241233
rect 147126 241159 147182 241168
rect 148336 225622 148364 256838
rect 148324 225616 148376 225622
rect 148324 225558 148376 225564
rect 147036 213376 147088 213382
rect 147036 213318 147088 213324
rect 146944 203856 146996 203862
rect 146944 203798 146996 203804
rect 144368 196920 144420 196926
rect 144368 196862 144420 196868
rect 144276 193928 144328 193934
rect 144276 193870 144328 193876
rect 142802 188456 142858 188465
rect 142802 188391 142858 188400
rect 141424 185768 141476 185774
rect 141424 185710 141476 185716
rect 148428 185706 148456 298250
rect 148508 296880 148560 296886
rect 148508 296822 148560 296828
rect 148520 191282 148548 296822
rect 148600 274780 148652 274786
rect 148600 274722 148652 274728
rect 148612 233102 148640 274722
rect 149716 238678 149744 391954
rect 151832 376689 151860 405062
rect 153108 396908 153160 396914
rect 153108 396850 153160 396856
rect 151818 376680 151874 376689
rect 151818 376615 151874 376624
rect 152554 376680 152610 376689
rect 152554 376615 152610 376624
rect 152568 375465 152596 376615
rect 152554 375456 152610 375465
rect 152554 375391 152610 375400
rect 152464 365832 152516 365838
rect 152464 365774 152516 365780
rect 151084 300892 151136 300898
rect 151084 300834 151136 300840
rect 149980 295452 150032 295458
rect 149980 295394 150032 295400
rect 149796 295384 149848 295390
rect 149796 295326 149848 295332
rect 149704 238672 149756 238678
rect 149704 238614 149756 238620
rect 148600 233096 148652 233102
rect 148600 233038 148652 233044
rect 148508 191276 148560 191282
rect 148508 191218 148560 191224
rect 148416 185700 148468 185706
rect 148416 185642 148468 185648
rect 149808 184482 149836 295326
rect 149888 289944 149940 289950
rect 149888 289886 149940 289892
rect 149900 194041 149928 289886
rect 149992 206582 150020 295394
rect 149980 206576 150032 206582
rect 149980 206518 150032 206524
rect 149886 194032 149942 194041
rect 149886 193967 149942 193976
rect 151096 186969 151124 300834
rect 151176 296744 151228 296750
rect 151176 296686 151228 296692
rect 151082 186960 151138 186969
rect 151082 186895 151138 186904
rect 149796 184476 149848 184482
rect 149796 184418 149848 184424
rect 151188 182889 151216 296686
rect 151268 254040 151320 254046
rect 151268 253982 151320 253988
rect 151280 235346 151308 253982
rect 152476 237250 152504 365774
rect 152568 349858 152596 375391
rect 152556 349852 152608 349858
rect 152556 349794 152608 349800
rect 152556 281648 152608 281654
rect 152556 281590 152608 281596
rect 152464 237244 152516 237250
rect 152464 237186 152516 237192
rect 151268 235340 151320 235346
rect 151268 235282 151320 235288
rect 151174 182880 151230 182889
rect 151174 182815 151230 182824
rect 138756 178696 138808 178702
rect 138756 178638 138808 178644
rect 148232 178152 148284 178158
rect 148232 178094 148284 178100
rect 134524 177948 134576 177954
rect 134524 177890 134576 177896
rect 132406 177576 132462 177585
rect 132406 177511 132462 177520
rect 133602 177576 133658 177585
rect 133602 177511 133658 177520
rect 134432 177064 134484 177070
rect 134432 177006 134484 177012
rect 134444 176769 134472 177006
rect 148244 176769 148272 178094
rect 112442 176760 112498 176769
rect 112442 176695 112498 176704
rect 125782 176760 125838 176769
rect 125782 176695 125838 176704
rect 127070 176760 127126 176769
rect 127070 176695 127126 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 130750 176760 130806 176769
rect 130750 176695 130806 176704
rect 134430 176760 134486 176769
rect 134430 176695 134486 176704
rect 135718 176760 135774 176769
rect 135718 176695 135720 176704
rect 135772 176695 135774 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 135720 176666 135772 176672
rect 129464 176316 129516 176322
rect 129464 176258 129516 176264
rect 119436 176248 119488 176254
rect 119436 176190 119488 176196
rect 115756 176180 115808 176186
rect 115756 176122 115808 176128
rect 111064 175976 111116 175982
rect 111064 175918 111116 175924
rect 98366 175400 98422 175409
rect 98366 175335 98422 175344
rect 100758 175400 100814 175409
rect 100758 175335 100814 175344
rect 115768 175001 115796 176122
rect 116952 175976 117004 175982
rect 116952 175918 117004 175924
rect 116964 175409 116992 175918
rect 116950 175400 117006 175409
rect 116950 175335 117006 175344
rect 119448 175001 119476 176190
rect 129476 175409 129504 176258
rect 152568 175953 152596 281590
rect 152648 245676 152700 245682
rect 152648 245618 152700 245624
rect 152660 191049 152688 245618
rect 153120 227662 153148 396850
rect 153844 391264 153896 391270
rect 153844 391206 153896 391212
rect 153856 244254 153884 391206
rect 155868 357740 155920 357746
rect 155868 357682 155920 357688
rect 153936 307828 153988 307834
rect 153936 307770 153988 307776
rect 153844 244248 153896 244254
rect 153844 244190 153896 244196
rect 153844 240168 153896 240174
rect 153844 240110 153896 240116
rect 153108 227656 153160 227662
rect 153108 227598 153160 227604
rect 153120 227050 153148 227598
rect 153108 227044 153160 227050
rect 153108 226986 153160 226992
rect 152646 191040 152702 191049
rect 152646 190975 152702 190984
rect 153856 189990 153884 240110
rect 153948 200802 153976 307770
rect 155316 299736 155368 299742
rect 155316 299678 155368 299684
rect 155224 287088 155276 287094
rect 155224 287030 155276 287036
rect 154028 269204 154080 269210
rect 154028 269146 154080 269152
rect 154040 214878 154068 269146
rect 154488 231192 154540 231198
rect 154488 231134 154540 231140
rect 154500 230450 154528 231134
rect 154488 230444 154540 230450
rect 154488 230386 154540 230392
rect 155236 229022 155264 287030
rect 155328 241466 155356 299678
rect 155316 241460 155368 241466
rect 155316 241402 155368 241408
rect 155224 229016 155276 229022
rect 155224 228958 155276 228964
rect 154028 214872 154080 214878
rect 154028 214814 154080 214820
rect 153936 200796 153988 200802
rect 153936 200738 153988 200744
rect 153844 189984 153896 189990
rect 153844 189926 153896 189932
rect 155880 184550 155908 357682
rect 155972 242282 156000 405062
rect 158732 401674 158760 405076
rect 159362 403608 159418 403617
rect 159362 403543 159418 403552
rect 158076 401668 158128 401674
rect 158076 401610 158128 401616
rect 158720 401668 158772 401674
rect 158720 401610 158772 401616
rect 156604 399560 156656 399566
rect 156604 399502 156656 399508
rect 156616 284986 156644 399502
rect 157984 396840 158036 396846
rect 157984 396782 158036 396788
rect 157248 329860 157300 329866
rect 157248 329802 157300 329808
rect 157156 303748 157208 303754
rect 157156 303690 157208 303696
rect 156604 284980 156656 284986
rect 156604 284922 156656 284928
rect 156604 256828 156656 256834
rect 156604 256770 156656 256776
rect 155960 242276 156012 242282
rect 155960 242218 156012 242224
rect 156616 239970 156644 256770
rect 156604 239964 156656 239970
rect 156604 239906 156656 239912
rect 157168 187270 157196 303690
rect 157156 187264 157208 187270
rect 157156 187206 157208 187212
rect 155868 184544 155920 184550
rect 155868 184486 155920 184492
rect 157260 183054 157288 329802
rect 157996 296857 158024 396782
rect 158088 364410 158116 401610
rect 158076 364404 158128 364410
rect 158076 364346 158128 364352
rect 158088 318102 158116 364346
rect 158628 345772 158680 345778
rect 158628 345714 158680 345720
rect 158076 318096 158128 318102
rect 158076 318038 158128 318044
rect 157982 296848 158038 296857
rect 157982 296783 158038 296792
rect 157996 296714 158024 296783
rect 157996 296686 158208 296714
rect 157984 292800 158036 292806
rect 157984 292742 158036 292748
rect 157996 199646 158024 292742
rect 158076 273284 158128 273290
rect 158076 273226 158128 273232
rect 158088 207874 158116 273226
rect 158180 237114 158208 296686
rect 158640 238649 158668 345714
rect 159376 264246 159404 403543
rect 161952 402830 161980 405076
rect 164252 405062 165186 405090
rect 161940 402824 161992 402830
rect 161940 402766 161992 402772
rect 162768 402824 162820 402830
rect 162768 402766 162820 402772
rect 162780 388278 162808 402766
rect 164148 402348 164200 402354
rect 164148 402290 164200 402296
rect 162124 388272 162176 388278
rect 162124 388214 162176 388220
rect 162768 388272 162820 388278
rect 162768 388214 162820 388220
rect 160836 374672 160888 374678
rect 160836 374614 160888 374620
rect 160744 364404 160796 364410
rect 160744 364346 160796 364352
rect 160756 363798 160784 364346
rect 160744 363792 160796 363798
rect 160744 363734 160796 363740
rect 160008 357672 160060 357678
rect 160008 357614 160060 357620
rect 159456 299668 159508 299674
rect 159456 299610 159508 299616
rect 159364 264240 159416 264246
rect 159364 264182 159416 264188
rect 158626 238640 158682 238649
rect 158626 238575 158682 238584
rect 158640 237425 158668 238575
rect 158626 237416 158682 237425
rect 158626 237351 158682 237360
rect 159376 237182 159404 264182
rect 159364 237176 159416 237182
rect 159364 237118 159416 237124
rect 158168 237108 158220 237114
rect 158168 237050 158220 237056
rect 159468 228410 159496 299610
rect 159456 228404 159508 228410
rect 159456 228346 159508 228352
rect 158168 227112 158220 227118
rect 158168 227054 158220 227060
rect 158076 207868 158128 207874
rect 158076 207810 158128 207816
rect 158180 200938 158208 227054
rect 158168 200932 158220 200938
rect 158168 200874 158220 200880
rect 157984 199640 158036 199646
rect 157984 199582 158036 199588
rect 160020 190058 160048 357614
rect 160744 340944 160796 340950
rect 160744 340886 160796 340892
rect 160100 280832 160152 280838
rect 160100 280774 160152 280780
rect 160112 278118 160140 280774
rect 160100 278112 160152 278118
rect 160100 278054 160152 278060
rect 160756 239426 160784 340886
rect 160848 299606 160876 374614
rect 161754 358048 161810 358057
rect 161754 357983 161810 357992
rect 161768 357513 161796 357983
rect 161478 357504 161534 357513
rect 161478 357439 161534 357448
rect 161754 357504 161810 357513
rect 161754 357439 161810 357448
rect 160836 299600 160888 299606
rect 160836 299542 160888 299548
rect 160848 284306 160876 299542
rect 160836 284300 160888 284306
rect 160836 284242 160888 284248
rect 161388 278112 161440 278118
rect 161388 278054 161440 278060
rect 160836 269136 160888 269142
rect 160836 269078 160888 269084
rect 160744 239420 160796 239426
rect 160744 239362 160796 239368
rect 160742 237416 160798 237425
rect 160742 237351 160798 237360
rect 160756 195294 160784 237351
rect 160848 198218 160876 269078
rect 160928 259480 160980 259486
rect 160928 259422 160980 259428
rect 160940 234054 160968 259422
rect 160928 234048 160980 234054
rect 160928 233990 160980 233996
rect 161400 229770 161428 278054
rect 161492 260846 161520 357439
rect 162136 319462 162164 388214
rect 162780 387870 162808 388214
rect 162768 387864 162820 387870
rect 162768 387806 162820 387812
rect 162216 363724 162268 363730
rect 162216 363666 162268 363672
rect 162228 329118 162256 363666
rect 163504 359508 163556 359514
rect 163504 359450 163556 359456
rect 162216 329112 162268 329118
rect 162216 329054 162268 329060
rect 162124 319456 162176 319462
rect 162124 319398 162176 319404
rect 162768 315308 162820 315314
rect 162768 315250 162820 315256
rect 162780 314809 162808 315250
rect 162766 314800 162822 314809
rect 162766 314735 162822 314744
rect 162124 302388 162176 302394
rect 162124 302330 162176 302336
rect 161480 260840 161532 260846
rect 161480 260782 161532 260788
rect 161480 229832 161532 229838
rect 161480 229774 161532 229780
rect 161388 229764 161440 229770
rect 161388 229706 161440 229712
rect 161492 224233 161520 229774
rect 161478 224224 161534 224233
rect 161478 224159 161534 224168
rect 160836 198212 160888 198218
rect 160836 198154 160888 198160
rect 160744 195288 160796 195294
rect 160744 195230 160796 195236
rect 160008 190052 160060 190058
rect 160008 189994 160060 190000
rect 157248 183048 157300 183054
rect 157248 182990 157300 182996
rect 162136 178673 162164 302330
rect 162214 298752 162270 298761
rect 162214 298687 162270 298696
rect 162228 182986 162256 298687
rect 162308 258120 162360 258126
rect 162308 258062 162360 258068
rect 162320 238678 162348 258062
rect 162400 255332 162452 255338
rect 162400 255274 162452 255280
rect 162308 238672 162360 238678
rect 162308 238614 162360 238620
rect 162412 237250 162440 255274
rect 163516 237289 163544 359450
rect 163596 334008 163648 334014
rect 163596 333950 163648 333956
rect 163608 321570 163636 333950
rect 163596 321564 163648 321570
rect 163596 321506 163648 321512
rect 163596 291848 163648 291854
rect 163596 291790 163648 291796
rect 163608 240106 163636 291790
rect 163596 240100 163648 240106
rect 163596 240042 163648 240048
rect 163502 237280 163558 237289
rect 162400 237244 162452 237250
rect 163502 237215 163558 237224
rect 162400 237186 162452 237192
rect 163516 227662 163544 237215
rect 163504 227656 163556 227662
rect 163504 227598 163556 227604
rect 163504 218952 163556 218958
rect 163504 218894 163556 218900
rect 162308 216096 162360 216102
rect 162308 216038 162360 216044
rect 162320 192545 162348 216038
rect 163516 195362 163544 218894
rect 164160 215286 164188 402290
rect 164252 372638 164280 405062
rect 165528 405000 165580 405006
rect 165528 404942 165580 404948
rect 164240 372632 164292 372638
rect 164240 372574 164292 372580
rect 164884 372632 164936 372638
rect 164884 372574 164936 372580
rect 164238 353424 164294 353433
rect 164238 353359 164294 353368
rect 164252 245614 164280 353359
rect 164896 322250 164924 372574
rect 165436 355020 165488 355026
rect 165436 354962 165488 354968
rect 165448 354657 165476 354962
rect 165434 354648 165490 354657
rect 165434 354583 165490 354592
rect 165448 353433 165476 354583
rect 165434 353424 165490 353433
rect 165434 353359 165490 353368
rect 164884 322244 164936 322250
rect 164884 322186 164936 322192
rect 164976 274712 165028 274718
rect 164976 274654 165028 274660
rect 164240 245608 164292 245614
rect 164240 245550 164292 245556
rect 164884 244996 164936 245002
rect 164884 244938 164936 244944
rect 164148 215280 164200 215286
rect 164148 215222 164200 215228
rect 164160 214742 164188 215222
rect 164148 214736 164200 214742
rect 164148 214678 164200 214684
rect 163504 195356 163556 195362
rect 163504 195298 163556 195304
rect 162400 194064 162452 194070
rect 162400 194006 162452 194012
rect 162306 192536 162362 192545
rect 162306 192471 162362 192480
rect 162216 182980 162268 182986
rect 162216 182922 162268 182928
rect 162122 178664 162178 178673
rect 162122 178599 162178 178608
rect 159916 178084 159968 178090
rect 159916 178026 159968 178032
rect 159928 176769 159956 178026
rect 159914 176760 159970 176769
rect 159914 176695 159970 176704
rect 162412 176633 162440 194006
rect 164896 181529 164924 244938
rect 164988 218958 165016 274654
rect 165540 241505 165568 404942
rect 168288 402280 168340 402286
rect 168288 402222 168340 402228
rect 166264 392692 166316 392698
rect 166264 392634 166316 392640
rect 166276 253910 166304 392634
rect 166816 377460 166868 377466
rect 166816 377402 166868 377408
rect 166828 282878 166856 377402
rect 168196 370592 168248 370598
rect 168196 370534 168248 370540
rect 166908 359032 166960 359038
rect 166908 358974 166960 358980
rect 166816 282872 166868 282878
rect 166816 282814 166868 282820
rect 166356 266416 166408 266422
rect 166356 266358 166408 266364
rect 166264 253904 166316 253910
rect 166264 253846 166316 253852
rect 165526 241496 165582 241505
rect 165526 241431 165582 241440
rect 165540 240825 165568 241431
rect 165526 240816 165582 240825
rect 165526 240751 165582 240760
rect 166368 234462 166396 266358
rect 166724 252612 166776 252618
rect 166724 252554 166776 252560
rect 166736 235414 166764 252554
rect 166816 249824 166868 249830
rect 166816 249766 166868 249772
rect 166724 235408 166776 235414
rect 166724 235350 166776 235356
rect 166356 234456 166408 234462
rect 166356 234398 166408 234404
rect 164976 218952 165028 218958
rect 164976 218894 165028 218900
rect 164882 181520 164938 181529
rect 164882 181455 164938 181464
rect 164332 180940 164384 180946
rect 164332 180882 164384 180888
rect 162398 176624 162454 176633
rect 162398 176559 162454 176568
rect 152554 175944 152610 175953
rect 152554 175879 152610 175888
rect 129462 175400 129518 175409
rect 129462 175335 129518 175344
rect 164344 175166 164372 180882
rect 166356 179648 166408 179654
rect 166356 179590 166408 179596
rect 165528 178220 165580 178226
rect 165528 178162 165580 178168
rect 165252 177064 165304 177070
rect 165252 177006 165304 177012
rect 165264 175234 165292 177006
rect 165252 175228 165304 175234
rect 165252 175170 165304 175176
rect 164332 175160 164384 175166
rect 164332 175102 164384 175108
rect 115754 174992 115810 175001
rect 115754 174927 115810 174936
rect 119434 174992 119490 175001
rect 119434 174927 119490 174936
rect 67546 129296 67602 129305
rect 67546 129231 67602 129240
rect 66166 128072 66222 128081
rect 66166 128007 66222 128016
rect 66180 127129 66208 128007
rect 64786 127120 64842 127129
rect 64786 127055 64842 127064
rect 66166 127120 66222 127129
rect 66166 127055 66222 127064
rect 63408 125656 63460 125662
rect 63408 125598 63460 125604
rect 63316 121508 63368 121514
rect 63316 121450 63368 121456
rect 63328 93770 63356 121450
rect 63316 93764 63368 93770
rect 63316 93706 63368 93712
rect 63420 86970 63448 125598
rect 64694 102232 64750 102241
rect 64694 102167 64750 102176
rect 63408 86964 63460 86970
rect 63408 86906 63460 86912
rect 64708 84182 64736 102167
rect 64800 93702 64828 127055
rect 66166 126304 66222 126313
rect 66166 126239 66222 126248
rect 66180 125662 66208 126239
rect 66168 125656 66220 125662
rect 66168 125598 66220 125604
rect 66166 125216 66222 125225
rect 66166 125151 66222 125160
rect 66074 122632 66130 122641
rect 66074 122567 66130 122576
rect 66088 121514 66116 122567
rect 66076 121508 66128 121514
rect 66076 121450 66128 121456
rect 64788 93696 64840 93702
rect 64788 93638 64840 93644
rect 66180 90982 66208 125151
rect 67454 123584 67510 123593
rect 67454 123519 67510 123528
rect 67362 120864 67418 120873
rect 67362 120799 67418 120808
rect 67376 91050 67404 120799
rect 67364 91044 67416 91050
rect 67364 90986 67416 90992
rect 66168 90976 66220 90982
rect 66168 90918 66220 90924
rect 67468 89729 67496 123519
rect 67560 94897 67588 129231
rect 67638 100736 67694 100745
rect 67638 100671 67694 100680
rect 67546 94888 67602 94897
rect 67546 94823 67602 94832
rect 67454 89720 67510 89729
rect 67454 89655 67510 89664
rect 67652 85542 67680 100671
rect 165540 173874 165568 178162
rect 166172 176316 166224 176322
rect 166172 176258 166224 176264
rect 165528 173868 165580 173874
rect 165528 173810 165580 173816
rect 166184 172514 166212 176258
rect 166264 176180 166316 176186
rect 166264 176122 166316 176128
rect 166172 172508 166224 172514
rect 166172 172450 166224 172456
rect 166276 165578 166304 176122
rect 166368 169726 166396 179590
rect 166828 177342 166856 249766
rect 166816 177336 166868 177342
rect 166920 177313 166948 358974
rect 167736 313268 167788 313274
rect 167736 313210 167788 313216
rect 167644 302252 167696 302258
rect 167644 302194 167696 302200
rect 167000 299464 167052 299470
rect 167000 299406 167052 299412
rect 167012 298790 167040 299406
rect 167000 298784 167052 298790
rect 167000 298726 167052 298732
rect 167000 291168 167052 291174
rect 167000 291110 167052 291116
rect 167012 290465 167040 291110
rect 166998 290456 167054 290465
rect 166998 290391 167054 290400
rect 167656 180198 167684 302194
rect 167748 301510 167776 313210
rect 167736 301504 167788 301510
rect 167736 301446 167788 301452
rect 167826 294264 167882 294273
rect 167826 294199 167882 294208
rect 167736 262268 167788 262274
rect 167736 262210 167788 262216
rect 167748 181558 167776 262210
rect 167840 238785 167868 294199
rect 168208 291174 168236 370534
rect 168300 299470 168328 402222
rect 168392 396982 168420 405076
rect 171048 405068 171100 405074
rect 171048 405010 171100 405016
rect 170956 398132 171008 398138
rect 170956 398074 171008 398080
rect 168380 396976 168432 396982
rect 168380 396918 168432 396924
rect 169116 367804 169168 367810
rect 169116 367746 169168 367752
rect 169024 316056 169076 316062
rect 169024 315998 169076 316004
rect 168288 299464 168340 299470
rect 168288 299406 168340 299412
rect 168196 291168 168248 291174
rect 168196 291110 168248 291116
rect 167920 285728 167972 285734
rect 167920 285670 167972 285676
rect 167826 238776 167882 238785
rect 167826 238711 167882 238720
rect 167932 232966 167960 285670
rect 168012 239420 168064 239426
rect 168012 239362 168064 239368
rect 167920 232960 167972 232966
rect 167920 232902 167972 232908
rect 168024 206514 168052 239362
rect 168012 206508 168064 206514
rect 168012 206450 168064 206456
rect 167920 186448 167972 186454
rect 167920 186390 167972 186396
rect 167828 182232 167880 182238
rect 167828 182174 167880 182180
rect 167736 181552 167788 181558
rect 167736 181494 167788 181500
rect 167644 180192 167696 180198
rect 167644 180134 167696 180140
rect 167736 179580 167788 179586
rect 167736 179522 167788 179528
rect 167644 178084 167696 178090
rect 167644 178026 167696 178032
rect 166816 177278 166868 177284
rect 166906 177304 166962 177313
rect 166906 177239 166962 177248
rect 166538 176624 166594 176633
rect 166538 176559 166594 176568
rect 166448 176248 166500 176254
rect 166448 176190 166500 176196
rect 166356 169720 166408 169726
rect 166356 169662 166408 169668
rect 166460 167006 166488 176190
rect 166552 175302 166580 176559
rect 166540 175296 166592 175302
rect 166540 175238 166592 175244
rect 166448 167000 166500 167006
rect 166448 166942 166500 166948
rect 166264 165572 166316 165578
rect 166264 165514 166316 165520
rect 167656 149054 167684 178026
rect 167748 168366 167776 179522
rect 167736 168360 167788 168366
rect 167736 168302 167788 168308
rect 167840 166938 167868 182174
rect 167932 173806 167960 186390
rect 169036 179314 169064 315998
rect 169128 292913 169156 367746
rect 170404 354884 170456 354890
rect 170404 354826 170456 354832
rect 169114 292904 169170 292913
rect 169114 292839 169170 292848
rect 169128 280158 169156 292839
rect 169298 292768 169354 292777
rect 169298 292703 169354 292712
rect 169116 280152 169168 280158
rect 169116 280094 169168 280100
rect 169208 278044 169260 278050
rect 169208 277986 169260 277992
rect 169220 233918 169248 277986
rect 169312 238542 169340 292703
rect 170416 288386 170444 354826
rect 170864 352708 170916 352714
rect 170864 352650 170916 352656
rect 170404 288380 170456 288386
rect 170404 288322 170456 288328
rect 169392 285796 169444 285802
rect 169392 285738 169444 285744
rect 169300 238536 169352 238542
rect 169300 238478 169352 238484
rect 169208 233912 169260 233918
rect 169208 233854 169260 233860
rect 169404 189854 169432 285738
rect 170404 281580 170456 281586
rect 170404 281522 170456 281528
rect 169760 231668 169812 231674
rect 169760 231610 169812 231616
rect 169772 231198 169800 231610
rect 169760 231192 169812 231198
rect 169760 231134 169812 231140
rect 170416 221542 170444 281522
rect 170770 231840 170826 231849
rect 170770 231775 170826 231784
rect 170404 221536 170456 221542
rect 170404 221478 170456 221484
rect 169760 208344 169812 208350
rect 169760 208286 169812 208292
rect 169772 207942 169800 208286
rect 169760 207936 169812 207942
rect 169760 207878 169812 207884
rect 169392 189848 169444 189854
rect 169392 189790 169444 189796
rect 169208 189168 169260 189174
rect 169208 189110 169260 189116
rect 169024 179308 169076 179314
rect 169024 179250 169076 179256
rect 169024 176112 169076 176118
rect 169024 176054 169076 176060
rect 167920 173800 167972 173806
rect 167920 173742 167972 173748
rect 167918 171592 167974 171601
rect 167918 171527 167974 171536
rect 167828 166932 167880 166938
rect 167828 166874 167880 166880
rect 167932 160818 167960 171527
rect 167920 160812 167972 160818
rect 167920 160754 167972 160760
rect 169036 155922 169064 176054
rect 169116 175976 169168 175982
rect 169116 175918 169168 175924
rect 169128 166870 169156 175918
rect 169116 166864 169168 166870
rect 169116 166806 169168 166812
rect 169220 160070 169248 189110
rect 170404 185020 170456 185026
rect 170404 184962 170456 184968
rect 169300 176792 169352 176798
rect 169300 176734 169352 176740
rect 169312 170406 169340 176734
rect 169300 170400 169352 170406
rect 169300 170342 169352 170348
rect 169208 160064 169260 160070
rect 169208 160006 169260 160012
rect 170416 157350 170444 184962
rect 170496 176860 170548 176866
rect 170496 176802 170548 176808
rect 170508 169046 170536 176802
rect 170496 169040 170548 169046
rect 170496 168982 170548 168988
rect 170404 157344 170456 157350
rect 170404 157286 170456 157292
rect 169024 155916 169076 155922
rect 169024 155858 169076 155864
rect 167644 149048 167696 149054
rect 167644 148990 167696 148996
rect 170404 144968 170456 144974
rect 170404 144910 170456 144916
rect 167644 143608 167696 143614
rect 167644 143550 167696 143556
rect 166264 133952 166316 133958
rect 166264 133894 166316 133900
rect 164884 99408 164936 99414
rect 164884 99350 164936 99356
rect 109038 94752 109094 94761
rect 109038 94687 109094 94696
rect 113730 94752 113786 94761
rect 113730 94687 113786 94696
rect 131946 94752 132002 94761
rect 131946 94687 132002 94696
rect 151726 94752 151782 94761
rect 151726 94687 151782 94696
rect 151910 94752 151966 94761
rect 151910 94687 151966 94696
rect 109052 93974 109080 94687
rect 109040 93968 109092 93974
rect 109040 93910 109092 93916
rect 113744 93906 113772 94687
rect 131960 94178 131988 94687
rect 131948 94172 132000 94178
rect 131948 94114 132000 94120
rect 151740 94042 151768 94687
rect 151924 94110 151952 94687
rect 151912 94104 151964 94110
rect 151912 94046 151964 94052
rect 151728 94036 151780 94042
rect 151728 93978 151780 93984
rect 113732 93900 113784 93906
rect 113732 93842 113784 93848
rect 121734 93664 121790 93673
rect 121734 93599 121790 93608
rect 102046 93528 102102 93537
rect 102046 93463 102102 93472
rect 107750 93528 107806 93537
rect 107750 93463 107806 93472
rect 102060 93158 102088 93463
rect 107764 93226 107792 93463
rect 121748 93362 121776 93599
rect 124494 93528 124550 93537
rect 124494 93463 124550 93472
rect 121736 93356 121788 93362
rect 121736 93298 121788 93304
rect 124508 93294 124536 93463
rect 124496 93288 124548 93294
rect 110142 93256 110198 93265
rect 107752 93220 107804 93226
rect 110142 93191 110198 93200
rect 119342 93256 119398 93265
rect 124496 93230 124548 93236
rect 119342 93191 119398 93200
rect 107752 93162 107804 93168
rect 102048 93152 102100 93158
rect 102048 93094 102100 93100
rect 74814 92440 74870 92449
rect 74814 92375 74870 92384
rect 85946 92440 86002 92449
rect 85946 92375 86002 92384
rect 94226 92440 94282 92449
rect 94226 92375 94282 92384
rect 101862 92440 101918 92449
rect 101862 92375 101918 92384
rect 74828 91118 74856 92375
rect 85026 91216 85082 91225
rect 85960 91186 85988 92375
rect 89074 91760 89130 91769
rect 89074 91695 89130 91704
rect 86774 91216 86830 91225
rect 85026 91151 85082 91160
rect 85948 91180 86000 91186
rect 74816 91112 74868 91118
rect 74816 91054 74868 91060
rect 67640 85536 67692 85542
rect 67640 85478 67692 85484
rect 85040 85474 85068 91151
rect 86774 91151 86830 91160
rect 87418 91216 87474 91225
rect 87418 91151 87474 91160
rect 85948 91122 86000 91128
rect 85028 85468 85080 85474
rect 85028 85410 85080 85416
rect 64696 84176 64748 84182
rect 64696 84118 64748 84124
rect 86788 82618 86816 91151
rect 87432 88194 87460 91151
rect 89088 89690 89116 91695
rect 94240 91322 94268 92375
rect 99286 91488 99342 91497
rect 99286 91423 99342 91432
rect 97906 91352 97962 91361
rect 94228 91316 94280 91322
rect 97906 91287 97962 91296
rect 99102 91352 99158 91361
rect 99102 91287 99158 91296
rect 94228 91258 94280 91264
rect 91006 91216 91062 91225
rect 91006 91151 91062 91160
rect 92386 91216 92442 91225
rect 92386 91151 92442 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 95054 91216 95110 91225
rect 95054 91151 95110 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97814 91216 97870 91225
rect 97814 91151 97870 91160
rect 89076 89684 89128 89690
rect 89076 89626 89128 89632
rect 91020 88330 91048 91151
rect 91008 88324 91060 88330
rect 91008 88266 91060 88272
rect 87420 88188 87472 88194
rect 87420 88130 87472 88136
rect 86776 82612 86828 82618
rect 86776 82554 86828 82560
rect 92400 81326 92428 91151
rect 92388 81320 92440 81326
rect 92388 81262 92440 81268
rect 80060 76560 80112 76566
rect 80060 76502 80112 76508
rect 64880 66904 64932 66910
rect 64880 66846 64932 66852
rect 58624 59356 58676 59362
rect 58624 59298 58676 59304
rect 63500 54528 63552 54534
rect 63500 54470 63552 54476
rect 60740 53100 60792 53106
rect 60740 53042 60792 53048
rect 59360 21480 59412 21486
rect 59360 21422 59412 21428
rect 53852 16546 54984 16574
rect 57992 16546 58480 16574
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3470
rect 54956 480 54984 16546
rect 56598 8936 56654 8945
rect 56598 8871 56654 8880
rect 56612 3602 56640 8871
rect 56600 3596 56652 3602
rect 56600 3538 56652 3544
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 56048 2100 56100 2106
rect 56048 2042 56100 2048
rect 56060 480 56088 2042
rect 57256 480 57284 3470
rect 58452 480 58480 16546
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59372 354 59400 21422
rect 60752 16574 60780 53042
rect 62120 24200 62172 24206
rect 62120 24142 62172 24148
rect 62132 16574 62160 24142
rect 63512 16574 63540 54470
rect 64892 16574 64920 66846
rect 69020 65544 69072 65550
rect 69020 65486 69072 65492
rect 67640 61396 67692 61402
rect 67640 61338 67692 61344
rect 60752 16546 60872 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 60844 480 60872 16546
rect 62028 7676 62080 7682
rect 62028 7618 62080 7624
rect 62040 480 62068 7618
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66720 14476 66772 14482
rect 66720 14418 66772 14424
rect 66732 480 66760 14418
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 61338
rect 69032 16574 69060 65486
rect 71780 64252 71832 64258
rect 71780 64194 71832 64200
rect 70400 55888 70452 55894
rect 70400 55830 70452 55836
rect 70412 16574 70440 55830
rect 71792 16574 71820 64194
rect 74540 57316 74592 57322
rect 74540 57258 74592 57264
rect 73160 29708 73212 29714
rect 73160 29650 73212 29656
rect 73172 16574 73200 29650
rect 74552 16574 74580 57258
rect 78680 36644 78732 36650
rect 78680 36586 78732 36592
rect 75920 31068 75972 31074
rect 75920 31010 75972 31016
rect 69032 16546 69152 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69124 480 69152 16546
rect 70308 6180 70360 6186
rect 70308 6122 70360 6128
rect 70320 480 70348 6122
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 31010
rect 77300 25560 77352 25566
rect 77300 25502 77352 25508
rect 77312 16574 77340 25502
rect 78692 16574 78720 36586
rect 80072 16574 80100 76502
rect 93780 75886 93808 91151
rect 95068 81258 95096 91151
rect 96540 85406 96568 91151
rect 96528 85400 96580 85406
rect 96528 85342 96580 85348
rect 95056 81252 95108 81258
rect 95056 81194 95108 81200
rect 97828 79830 97856 91151
rect 97816 79824 97868 79830
rect 97816 79766 97868 79772
rect 97920 78606 97948 91287
rect 99116 79762 99144 91287
rect 99194 91216 99250 91225
rect 99194 91151 99250 91160
rect 99104 79756 99156 79762
rect 99104 79698 99156 79704
rect 97908 78600 97960 78606
rect 99208 78577 99236 91151
rect 97908 78542 97960 78548
rect 99194 78568 99250 78577
rect 99194 78503 99250 78512
rect 99300 77246 99328 91423
rect 101876 91254 101904 92375
rect 104530 91624 104586 91633
rect 104530 91559 104586 91568
rect 106922 91624 106978 91633
rect 106922 91559 106978 91568
rect 101864 91248 101916 91254
rect 99930 91216 99986 91225
rect 99930 91151 99986 91160
rect 100666 91216 100722 91225
rect 101864 91190 101916 91196
rect 102046 91216 102102 91225
rect 100666 91151 100722 91160
rect 102046 91151 102102 91160
rect 102966 91216 103022 91225
rect 102966 91151 103022 91160
rect 103426 91216 103482 91225
rect 103426 91151 103482 91160
rect 99944 86902 99972 91151
rect 99932 86896 99984 86902
rect 99932 86838 99984 86844
rect 100680 82822 100708 91151
rect 100668 82816 100720 82822
rect 100668 82758 100720 82764
rect 102060 79966 102088 91151
rect 102980 86766 103008 91151
rect 102968 86760 103020 86766
rect 102968 86702 103020 86708
rect 103440 82550 103468 91151
rect 104544 89486 104572 91559
rect 104622 91216 104678 91225
rect 104622 91151 104678 91160
rect 106186 91216 106242 91225
rect 106186 91151 106242 91160
rect 106646 91216 106702 91225
rect 106646 91151 106702 91160
rect 104532 89480 104584 89486
rect 104532 89422 104584 89428
rect 104636 86873 104664 91151
rect 104622 86864 104678 86873
rect 104622 86799 104678 86808
rect 106200 83978 106228 91151
rect 106660 88262 106688 91151
rect 106936 89418 106964 91559
rect 106924 89412 106976 89418
rect 106924 89354 106976 89360
rect 106648 88256 106700 88262
rect 106648 88198 106700 88204
rect 110156 88126 110184 93191
rect 119356 92478 119384 93191
rect 119344 92472 119396 92478
rect 115202 92440 115258 92449
rect 115202 92375 115258 92384
rect 115478 92440 115534 92449
rect 119344 92414 119396 92420
rect 120354 92440 120410 92449
rect 115478 92375 115534 92384
rect 120354 92375 120356 92384
rect 112350 91760 112406 91769
rect 112350 91695 112406 91704
rect 110326 91216 110382 91225
rect 110326 91151 110382 91160
rect 110694 91216 110750 91225
rect 110694 91151 110750 91160
rect 111706 91216 111762 91225
rect 111706 91151 111762 91160
rect 110144 88120 110196 88126
rect 110144 88062 110196 88068
rect 110340 84153 110368 91151
rect 110708 88233 110736 91151
rect 110694 88224 110750 88233
rect 110694 88159 110750 88168
rect 110326 84144 110382 84153
rect 110326 84079 110382 84088
rect 106188 83972 106240 83978
rect 106188 83914 106240 83920
rect 103428 82544 103480 82550
rect 103428 82486 103480 82492
rect 102048 79960 102100 79966
rect 102048 79902 102100 79908
rect 99288 77240 99340 77246
rect 99288 77182 99340 77188
rect 93768 75880 93820 75886
rect 93768 75822 93820 75828
rect 111720 75818 111748 91151
rect 112364 89554 112392 91695
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 112444 91112 112496 91118
rect 112444 91054 112496 91060
rect 112352 89548 112404 89554
rect 112352 89490 112404 89496
rect 112456 84114 112484 91054
rect 112444 84108 112496 84114
rect 112444 84050 112496 84056
rect 114480 77178 114508 91151
rect 115216 90846 115244 92375
rect 115492 92342 115520 92375
rect 120408 92375 120410 92384
rect 124126 92440 124182 92449
rect 124126 92375 124182 92384
rect 125966 92440 126022 92449
rect 125966 92375 126022 92384
rect 133142 92440 133198 92449
rect 133142 92375 133198 92384
rect 151726 92440 151782 92449
rect 151726 92375 151782 92384
rect 120356 92346 120408 92352
rect 115480 92336 115532 92342
rect 115480 92278 115532 92284
rect 123942 91760 123998 91769
rect 123942 91695 123998 91704
rect 122838 91488 122894 91497
rect 122838 91423 122894 91432
rect 118238 91352 118294 91361
rect 118238 91287 118294 91296
rect 120724 91316 120776 91322
rect 115754 91216 115810 91225
rect 115754 91151 115810 91160
rect 116766 91216 116822 91225
rect 116766 91151 116822 91160
rect 117134 91216 117190 91225
rect 117134 91151 117190 91160
rect 115204 90840 115256 90846
rect 115204 90782 115256 90788
rect 115768 82686 115796 91151
rect 116780 85202 116808 91151
rect 117148 86834 117176 91151
rect 117136 86828 117188 86834
rect 117136 86770 117188 86776
rect 118252 85338 118280 91287
rect 120724 91258 120776 91264
rect 118606 91216 118662 91225
rect 118606 91151 118662 91160
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 118240 85332 118292 85338
rect 118240 85274 118292 85280
rect 116768 85196 116820 85202
rect 116768 85138 116820 85144
rect 115756 82680 115808 82686
rect 115756 82622 115808 82628
rect 118620 78470 118648 91151
rect 120000 84046 120028 91151
rect 119988 84040 120040 84046
rect 119988 83982 120040 83988
rect 120736 79898 120764 91258
rect 121090 91216 121146 91225
rect 120816 91180 120868 91186
rect 121090 91151 121146 91160
rect 122378 91216 122434 91225
rect 122378 91151 122434 91160
rect 120816 91122 120868 91128
rect 120828 81122 120856 91122
rect 121104 87990 121132 91151
rect 121092 87984 121144 87990
rect 121092 87926 121144 87932
rect 122392 86698 122420 91151
rect 122852 90778 122880 91423
rect 122840 90772 122892 90778
rect 122840 90714 122892 90720
rect 123956 89622 123984 91695
rect 124140 90914 124168 92375
rect 125980 92138 126008 92375
rect 133156 92274 133184 92375
rect 133144 92268 133196 92274
rect 133144 92210 133196 92216
rect 151740 92206 151768 92375
rect 151728 92200 151780 92206
rect 151728 92142 151780 92148
rect 125968 92132 126020 92138
rect 125968 92074 126020 92080
rect 151726 91760 151782 91769
rect 151726 91695 151782 91704
rect 126610 91624 126666 91633
rect 126610 91559 126666 91568
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 124128 90908 124180 90914
rect 124128 90850 124180 90856
rect 123944 89616 123996 89622
rect 123944 89558 123996 89564
rect 122380 86692 122432 86698
rect 122380 86634 122432 86640
rect 120816 81116 120868 81122
rect 120816 81058 120868 81064
rect 120724 79892 120776 79898
rect 120724 79834 120776 79840
rect 125520 78538 125548 91151
rect 126624 89350 126652 91559
rect 127624 91248 127676 91254
rect 126886 91216 126942 91225
rect 127624 91190 127676 91196
rect 129646 91216 129702 91225
rect 126886 91151 126942 91160
rect 126612 89344 126664 89350
rect 126612 89286 126664 89292
rect 126900 82754 126928 91151
rect 126888 82748 126940 82754
rect 126888 82690 126940 82696
rect 125508 78532 125560 78538
rect 125508 78474 125560 78480
rect 118608 78464 118660 78470
rect 118608 78406 118660 78412
rect 114468 77172 114520 77178
rect 114468 77114 114520 77120
rect 115940 76628 115992 76634
rect 115940 76570 115992 76576
rect 111708 75812 111760 75818
rect 111708 75754 111760 75760
rect 98000 75200 98052 75206
rect 98000 75142 98052 75148
rect 81440 73908 81492 73914
rect 81440 73850 81492 73856
rect 81452 16574 81480 73850
rect 85580 72548 85632 72554
rect 85580 72490 85632 72496
rect 82820 61464 82872 61470
rect 82820 61406 82872 61412
rect 82832 16574 82860 61406
rect 84200 50448 84252 50454
rect 84200 50390 84252 50396
rect 77312 16546 77432 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77404 480 77432 16546
rect 78128 10328 78180 10334
rect 78128 10270 78180 10276
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 10270
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 50390
rect 85592 6914 85620 72490
rect 88338 69592 88394 69601
rect 88338 69527 88394 69536
rect 85672 60036 85724 60042
rect 85672 59978 85724 59984
rect 85684 16574 85712 59978
rect 86960 28348 87012 28354
rect 86960 28290 87012 28296
rect 86972 16574 87000 28290
rect 88352 16574 88380 69527
rect 92480 68400 92532 68406
rect 92480 68342 92532 68348
rect 89720 58676 89772 58682
rect 89720 58618 89772 58624
rect 89732 16574 89760 58618
rect 91100 19984 91152 19990
rect 91100 19926 91152 19932
rect 91112 16574 91140 19926
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 68342
rect 93860 57248 93912 57254
rect 93860 57190 93912 57196
rect 93872 6914 93900 57190
rect 96620 55956 96672 55962
rect 96620 55898 96672 55904
rect 93952 32428 94004 32434
rect 93952 32370 94004 32376
rect 93964 16574 93992 32370
rect 95240 17332 95292 17338
rect 95240 17274 95292 17280
rect 95252 16574 95280 17274
rect 96632 16574 96660 55898
rect 98012 16574 98040 75142
rect 113180 71188 113232 71194
rect 113180 71130 113232 71136
rect 99380 66972 99432 66978
rect 99380 66914 99432 66920
rect 99392 16574 99420 66914
rect 106280 65612 106332 65618
rect 106280 65554 106332 65560
rect 100760 54596 100812 54602
rect 100760 54538 100812 54544
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 54538
rect 103520 53168 103572 53174
rect 103520 53110 103572 53116
rect 102140 49088 102192 49094
rect 102140 49030 102192 49036
rect 102152 3602 102180 49030
rect 102232 43512 102284 43518
rect 102232 43454 102284 43460
rect 102140 3596 102192 3602
rect 102140 3538 102192 3544
rect 102244 480 102272 43454
rect 103532 16574 103560 53110
rect 104900 31136 104952 31142
rect 104900 31078 104952 31084
rect 104912 16574 104940 31078
rect 106292 16574 106320 65554
rect 110420 62892 110472 62898
rect 110420 62834 110472 62840
rect 107660 51808 107712 51814
rect 107660 51750 107712 51756
rect 107672 16574 107700 51750
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103348 480 103376 3538
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109040 11824 109092 11830
rect 109040 11766 109092 11772
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 11766
rect 110432 6914 110460 62834
rect 110512 40792 110564 40798
rect 110512 40734 110564 40740
rect 110524 16574 110552 40734
rect 113192 16574 113220 71130
rect 114560 18624 114612 18630
rect 114560 18566 114612 18572
rect 114572 16574 114600 18566
rect 115952 16574 115980 76570
rect 127636 74526 127664 91190
rect 129646 91151 129702 91160
rect 131026 91216 131082 91225
rect 131026 91151 131082 91160
rect 135074 91216 135130 91225
rect 135074 91151 135130 91160
rect 135902 91216 135958 91225
rect 135902 91151 135958 91160
rect 129660 83910 129688 91151
rect 129648 83904 129700 83910
rect 129648 83846 129700 83852
rect 131040 81190 131068 91151
rect 135088 85270 135116 91151
rect 135916 88058 135944 91151
rect 151740 90710 151768 91695
rect 151728 90704 151780 90710
rect 151728 90646 151780 90652
rect 164896 88194 164924 99350
rect 166276 88233 166304 133894
rect 166356 125656 166408 125662
rect 166356 125598 166408 125604
rect 166368 89350 166396 125598
rect 166448 118720 166500 118726
rect 166448 118662 166500 118668
rect 166460 90846 166488 118662
rect 166540 98048 166592 98054
rect 166540 97990 166592 97996
rect 166448 90840 166500 90846
rect 166448 90782 166500 90788
rect 166356 89344 166408 89350
rect 166356 89286 166408 89292
rect 166262 88224 166318 88233
rect 164884 88188 164936 88194
rect 166262 88159 166318 88168
rect 164884 88130 164936 88136
rect 135904 88052 135956 88058
rect 135904 87994 135956 88000
rect 135076 85264 135128 85270
rect 135076 85206 135128 85212
rect 166552 82618 166580 97990
rect 167656 83910 167684 143550
rect 169116 136672 169168 136678
rect 169116 136614 169168 136620
rect 169024 135312 169076 135318
rect 169024 135254 169076 135260
rect 167736 124228 167788 124234
rect 167736 124170 167788 124176
rect 167748 90778 167776 124170
rect 167828 117360 167880 117366
rect 167828 117302 167880 117308
rect 167736 90772 167788 90778
rect 167736 90714 167788 90720
rect 167840 88126 167868 117302
rect 167920 111784 167972 111790
rect 167918 111752 167920 111761
rect 167972 111752 167974 111761
rect 167918 111687 167974 111696
rect 168104 110424 168156 110430
rect 168104 110366 168156 110372
rect 168116 110129 168144 110366
rect 168102 110120 168158 110129
rect 168102 110055 168158 110064
rect 168012 109064 168064 109070
rect 168012 109006 168064 109012
rect 167920 108996 167972 109002
rect 167920 108938 167972 108944
rect 167932 108769 167960 108938
rect 167918 108760 167974 108769
rect 167918 108695 167974 108704
rect 168024 103514 168052 109006
rect 167932 103486 168052 103514
rect 167828 88120 167880 88126
rect 167828 88062 167880 88068
rect 167932 85406 167960 103486
rect 167920 85400 167972 85406
rect 167920 85342 167972 85348
rect 167644 83904 167696 83910
rect 167644 83846 167696 83852
rect 166540 82612 166592 82618
rect 166540 82554 166592 82560
rect 131028 81184 131080 81190
rect 131028 81126 131080 81132
rect 169036 77178 169064 135254
rect 169128 85202 169156 136614
rect 169300 116068 169352 116074
rect 169300 116010 169352 116016
rect 169208 116000 169260 116006
rect 169208 115942 169260 115948
rect 169220 93226 169248 115942
rect 169312 93974 169340 116010
rect 170416 94178 170444 144910
rect 170496 122868 170548 122874
rect 170496 122810 170548 122816
rect 170404 94172 170456 94178
rect 170404 94114 170456 94120
rect 169300 93968 169352 93974
rect 169300 93910 169352 93916
rect 169208 93220 169260 93226
rect 169208 93162 169260 93168
rect 170508 87990 170536 122810
rect 170784 113830 170812 231775
rect 170876 207942 170904 352650
rect 170968 313274 170996 398074
rect 170956 313268 171008 313274
rect 170956 313210 171008 313216
rect 170956 257372 171008 257378
rect 170956 257314 171008 257320
rect 170864 207936 170916 207942
rect 170864 207878 170916 207884
rect 170772 113824 170824 113830
rect 170772 113766 170824 113772
rect 170588 113212 170640 113218
rect 170588 113154 170640 113160
rect 170600 89486 170628 113154
rect 170968 102814 170996 257314
rect 171060 231674 171088 405010
rect 171612 402354 171640 405076
rect 171600 402348 171652 402354
rect 171600 402290 171652 402296
rect 173716 400920 173768 400926
rect 173716 400862 173768 400868
rect 171968 366376 172020 366382
rect 171968 366318 172020 366324
rect 171784 361684 171836 361690
rect 171784 361626 171836 361632
rect 171796 345710 171824 361626
rect 171876 360256 171928 360262
rect 171876 360198 171928 360204
rect 171784 345704 171836 345710
rect 171784 345646 171836 345652
rect 171784 303680 171836 303686
rect 171784 303622 171836 303628
rect 171048 231668 171100 231674
rect 171048 231610 171100 231616
rect 171796 127634 171824 303622
rect 171888 295361 171916 360198
rect 171980 356318 172008 366318
rect 172060 358964 172112 358970
rect 172060 358906 172112 358912
rect 171968 356312 172020 356318
rect 171968 356254 172020 356260
rect 171874 295352 171930 295361
rect 171874 295287 171930 295296
rect 171980 262206 172008 356254
rect 172072 351218 172100 358906
rect 172060 351212 172112 351218
rect 172060 351154 172112 351160
rect 172426 295352 172482 295361
rect 172426 295287 172482 295296
rect 172152 289876 172204 289882
rect 172152 289818 172204 289824
rect 171968 262200 172020 262206
rect 171968 262142 172020 262148
rect 171968 258732 172020 258738
rect 171968 258674 172020 258680
rect 171980 233986 172008 258674
rect 172060 244928 172112 244934
rect 172060 244870 172112 244876
rect 171968 233980 172020 233986
rect 171968 233922 172020 233928
rect 172072 230450 172100 244870
rect 172060 230444 172112 230450
rect 172060 230386 172112 230392
rect 172164 179382 172192 289818
rect 172440 288386 172468 295287
rect 173728 294642 173756 400862
rect 173808 399628 173860 399634
rect 173808 399570 173860 399576
rect 173716 294636 173768 294642
rect 173716 294578 173768 294584
rect 173728 294001 173756 294578
rect 173714 293992 173770 294001
rect 173714 293927 173770 293936
rect 172428 288380 172480 288386
rect 172428 288322 172480 288328
rect 173256 282940 173308 282946
rect 173256 282882 173308 282888
rect 173164 279472 173216 279478
rect 173164 279414 173216 279420
rect 172334 255232 172390 255241
rect 172334 255167 172390 255176
rect 172348 253978 172376 255167
rect 172336 253972 172388 253978
rect 172336 253914 172388 253920
rect 173176 187134 173204 279414
rect 173268 231198 173296 282882
rect 173820 238610 173848 399570
rect 174832 399566 174860 405076
rect 178052 404462 178080 405076
rect 181286 405062 181484 405090
rect 178040 404456 178092 404462
rect 178040 404398 178092 404404
rect 176566 403744 176622 403753
rect 176566 403679 176622 403688
rect 174820 399560 174872 399566
rect 174820 399502 174872 399508
rect 175188 395412 175240 395418
rect 175188 395354 175240 395360
rect 174636 357468 174688 357474
rect 174636 357410 174688 357416
rect 174544 356244 174596 356250
rect 174544 356186 174596 356192
rect 174556 248402 174584 356186
rect 174648 304298 174676 357410
rect 175200 354414 175228 395354
rect 176476 392624 176528 392630
rect 176476 392566 176528 392572
rect 175188 354408 175240 354414
rect 175188 354350 175240 354356
rect 175200 352578 175228 354350
rect 175188 352572 175240 352578
rect 175188 352514 175240 352520
rect 175188 351960 175240 351966
rect 175188 351902 175240 351908
rect 175096 316464 175148 316470
rect 175096 316406 175148 316412
rect 174636 304292 174688 304298
rect 174636 304234 174688 304240
rect 174636 299532 174688 299538
rect 174636 299474 174688 299480
rect 174648 295322 174676 299474
rect 174636 295316 174688 295322
rect 174636 295258 174688 295264
rect 174636 292664 174688 292670
rect 174636 292606 174688 292612
rect 174544 248396 174596 248402
rect 174544 248338 174596 248344
rect 173808 238604 173860 238610
rect 173808 238546 173860 238552
rect 173820 237454 173848 238546
rect 174648 238474 174676 292606
rect 174636 238468 174688 238474
rect 174636 238410 174688 238416
rect 173808 237448 173860 237454
rect 173808 237390 173860 237396
rect 173256 231192 173308 231198
rect 173256 231134 173308 231140
rect 173164 187128 173216 187134
rect 173164 187070 173216 187076
rect 173256 186380 173308 186386
rect 173256 186322 173308 186328
rect 172152 179376 172204 179382
rect 172152 179318 172204 179324
rect 173164 176996 173216 177002
rect 173164 176938 173216 176944
rect 171876 176044 171928 176050
rect 171876 175986 171928 175992
rect 171888 157282 171916 175986
rect 173176 171086 173204 176938
rect 173164 171080 173216 171086
rect 173164 171022 173216 171028
rect 173268 160002 173296 186322
rect 173256 159996 173308 160002
rect 173256 159938 173308 159944
rect 171876 157276 171928 157282
rect 171876 157218 171928 157224
rect 172060 135380 172112 135386
rect 172060 135322 172112 135328
rect 171876 129804 171928 129810
rect 171876 129746 171928 129752
rect 171784 127628 171836 127634
rect 171784 127570 171836 127576
rect 171784 120760 171836 120766
rect 171784 120702 171836 120708
rect 170956 102808 171008 102814
rect 170956 102750 171008 102756
rect 170680 101448 170732 101454
rect 170680 101390 170732 101396
rect 170692 92342 170720 101390
rect 170680 92336 170732 92342
rect 170680 92278 170732 92284
rect 171796 92138 171824 120702
rect 171784 92132 171836 92138
rect 171784 92074 171836 92080
rect 170588 89480 170640 89486
rect 170588 89422 170640 89428
rect 170496 87984 170548 87990
rect 170496 87926 170548 87932
rect 169116 85196 169168 85202
rect 169116 85138 169168 85144
rect 171888 82550 171916 129746
rect 171968 127016 172020 127022
rect 171968 126958 172020 126964
rect 171876 82544 171928 82550
rect 171876 82486 171928 82492
rect 171980 79762 172008 126958
rect 172072 93945 172100 135322
rect 173164 132524 173216 132530
rect 173164 132466 173216 132472
rect 172058 93936 172114 93945
rect 172058 93871 172114 93880
rect 173176 89418 173204 132466
rect 174544 129872 174596 129878
rect 174544 129814 174596 129820
rect 173348 122120 173400 122126
rect 173348 122062 173400 122068
rect 173256 114572 173308 114578
rect 173256 114514 173308 114520
rect 173164 89412 173216 89418
rect 173164 89354 173216 89360
rect 173268 83978 173296 114514
rect 173360 92177 173388 122062
rect 173440 100768 173492 100774
rect 173440 100710 173492 100716
rect 173346 92168 173402 92177
rect 173346 92103 173402 92112
rect 173452 85474 173480 100710
rect 174556 93158 174584 129814
rect 174636 106344 174688 106350
rect 174636 106286 174688 106292
rect 174544 93152 174596 93158
rect 174544 93094 174596 93100
rect 173440 85468 173492 85474
rect 173440 85410 173492 85416
rect 173256 83972 173308 83978
rect 173256 83914 173308 83920
rect 171968 79756 172020 79762
rect 171968 79698 172020 79704
rect 169024 77172 169076 77178
rect 169024 77114 169076 77120
rect 174648 75886 174676 106286
rect 174636 75880 174688 75886
rect 174636 75822 174688 75828
rect 127624 74520 127676 74526
rect 127624 74462 127676 74468
rect 117320 62824 117372 62830
rect 117320 62766 117372 62772
rect 110524 16546 111656 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 112352 15904 112404 15910
rect 112352 15846 112404 15852
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 15846
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 62766
rect 120080 58744 120132 58750
rect 120080 58686 120132 58692
rect 118700 42152 118752 42158
rect 118700 42094 118752 42100
rect 118712 16574 118740 42094
rect 120092 16574 120120 58686
rect 124220 49020 124272 49026
rect 124220 48962 124272 48968
rect 124232 16574 124260 48962
rect 128360 35284 128412 35290
rect 128360 35226 128412 35232
rect 128372 16574 128400 35226
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 124232 16546 124720 16574
rect 128372 16546 128952 16574
rect 118804 480 118832 16546
rect 119896 13116 119948 13122
rect 119896 13058 119948 13064
rect 119908 480 119936 13058
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122288 14544 122340 14550
rect 122288 14486 122340 14492
rect 122300 480 122328 14486
rect 123484 3596 123536 3602
rect 123484 3538 123536 3544
rect 123496 480 123524 3538
rect 124692 480 124720 16546
rect 125874 3360 125930 3369
rect 125874 3295 125930 3304
rect 125888 480 125916 3295
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 136456 6248 136508 6254
rect 136456 6190 136508 6196
rect 136468 480 136496 6190
rect 175108 4894 175136 316406
rect 175200 20058 175228 351902
rect 176488 333266 176516 392566
rect 176580 346338 176608 403679
rect 177856 400988 177908 400994
rect 177856 400930 177908 400936
rect 176660 354408 176712 354414
rect 176658 354376 176660 354385
rect 176712 354376 176714 354385
rect 176658 354311 176714 354320
rect 177578 352200 177634 352209
rect 177578 352135 177634 352144
rect 177592 351966 177620 352135
rect 177580 351960 177632 351966
rect 177580 351902 177632 351908
rect 176658 348120 176714 348129
rect 176658 348055 176714 348064
rect 176672 347818 176700 348055
rect 176660 347812 176712 347818
rect 176660 347754 176712 347760
rect 176580 346310 176700 346338
rect 176672 345778 176700 346310
rect 176660 345772 176712 345778
rect 176660 345714 176712 345720
rect 176672 345545 176700 345714
rect 176658 345536 176714 345545
rect 176658 345471 176714 345480
rect 176566 336560 176622 336569
rect 176566 336495 176622 336504
rect 176476 333260 176528 333266
rect 176476 333202 176528 333208
rect 176488 332625 176516 333202
rect 176474 332616 176530 332625
rect 176474 332551 176530 332560
rect 176474 323640 176530 323649
rect 176474 323575 176530 323584
rect 176016 292596 176068 292602
rect 176016 292538 176068 292544
rect 176028 238610 176056 292538
rect 176108 251252 176160 251258
rect 176108 251194 176160 251200
rect 176016 238604 176068 238610
rect 176016 238546 176068 238552
rect 175924 237448 175976 237454
rect 175924 237390 175976 237396
rect 175936 93838 175964 237390
rect 176120 235890 176148 251194
rect 176108 235884 176160 235890
rect 176108 235826 176160 235832
rect 176016 122936 176068 122942
rect 176016 122878 176068 122884
rect 175924 93832 175976 93838
rect 175924 93774 175976 93780
rect 176028 93362 176056 122878
rect 176016 93356 176068 93362
rect 176016 93298 176068 93304
rect 176488 83502 176516 323575
rect 176476 83496 176528 83502
rect 176476 83438 176528 83444
rect 176580 25634 176608 336495
rect 176658 334520 176714 334529
rect 176658 334455 176714 334464
rect 176672 334014 176700 334455
rect 176660 334008 176712 334014
rect 176660 333950 176712 333956
rect 176658 330440 176714 330449
rect 176658 330375 176714 330384
rect 176672 329866 176700 330375
rect 176660 329860 176712 329866
rect 176660 329802 176712 329808
rect 176660 327140 176712 327146
rect 176660 327082 176712 327088
rect 176672 325825 176700 327082
rect 176658 325816 176714 325825
rect 176658 325751 176714 325760
rect 177670 318880 177726 318889
rect 177670 318815 177726 318824
rect 177578 316840 177634 316849
rect 177578 316775 177634 316784
rect 177592 316470 177620 316775
rect 177580 316464 177632 316470
rect 177580 316406 177632 316412
rect 176660 315308 176712 315314
rect 176660 315250 176712 315256
rect 176672 314945 176700 315250
rect 176658 314936 176714 314945
rect 176658 314871 176714 314880
rect 176660 313268 176712 313274
rect 176660 313210 176712 313216
rect 176672 312905 176700 313210
rect 176658 312896 176714 312905
rect 176658 312831 176714 312840
rect 176658 310040 176714 310049
rect 176658 309975 176714 309984
rect 176672 309874 176700 309975
rect 176660 309868 176712 309874
rect 176660 309810 176712 309816
rect 176658 303920 176714 303929
rect 176658 303855 176714 303864
rect 176672 303754 176700 303855
rect 176660 303748 176712 303754
rect 176660 303690 176712 303696
rect 176660 299464 176712 299470
rect 176660 299406 176712 299412
rect 176672 299305 176700 299406
rect 176658 299296 176714 299305
rect 176658 299231 176714 299240
rect 176660 297492 176712 297498
rect 176660 297434 176712 297440
rect 176672 297265 176700 297434
rect 176658 297256 176714 297265
rect 176658 297191 176714 297200
rect 176660 295316 176712 295322
rect 176660 295258 176712 295264
rect 176672 295225 176700 295258
rect 176658 295216 176714 295225
rect 176658 295151 176714 295160
rect 176660 291168 176712 291174
rect 176660 291110 176712 291116
rect 176672 290465 176700 291110
rect 176658 290456 176714 290465
rect 176658 290391 176714 290400
rect 176658 288416 176714 288425
rect 176658 288351 176660 288360
rect 176712 288351 176714 288360
rect 176660 288322 176712 288328
rect 176660 284300 176712 284306
rect 176660 284242 176712 284248
rect 176672 283665 176700 284242
rect 176658 283656 176714 283665
rect 176658 283591 176714 283600
rect 176660 282872 176712 282878
rect 176660 282814 176712 282820
rect 176672 281625 176700 282814
rect 176658 281616 176714 281625
rect 176658 281551 176714 281560
rect 176752 280152 176804 280158
rect 176752 280094 176804 280100
rect 176764 279585 176792 280094
rect 176750 279576 176806 279585
rect 176750 279511 176806 279520
rect 176660 278112 176712 278118
rect 176660 278054 176712 278060
rect 176672 277545 176700 278054
rect 176658 277536 176714 277545
rect 176658 277471 176714 277480
rect 176660 276004 176712 276010
rect 176660 275946 176712 275952
rect 176672 274825 176700 275946
rect 176658 274816 176714 274825
rect 176658 274751 176714 274760
rect 176658 272640 176714 272649
rect 176658 272575 176714 272584
rect 176672 272542 176700 272575
rect 176660 272536 176712 272542
rect 176660 272478 176712 272484
rect 176660 262132 176712 262138
rect 176660 262074 176712 262080
rect 176672 261905 176700 262074
rect 176658 261896 176714 261905
rect 176658 261831 176714 261840
rect 176658 257000 176714 257009
rect 176658 256935 176714 256944
rect 176672 256766 176700 256935
rect 176660 256760 176712 256766
rect 176660 256702 176712 256708
rect 176658 254960 176714 254969
rect 176658 254895 176714 254904
rect 176672 253978 176700 254895
rect 176660 253972 176712 253978
rect 176660 253914 176712 253920
rect 176658 252920 176714 252929
rect 176658 252855 176714 252864
rect 176672 252618 176700 252855
rect 176660 252612 176712 252618
rect 176660 252554 176712 252560
rect 176658 250880 176714 250889
rect 176658 250815 176714 250824
rect 176672 249830 176700 250815
rect 176660 249824 176712 249830
rect 176660 249766 176712 249772
rect 176660 247036 176712 247042
rect 176660 246978 176712 246984
rect 176672 246265 176700 246978
rect 176658 246256 176714 246265
rect 176658 246191 176714 246200
rect 177684 225690 177712 318815
rect 177868 305969 177896 400930
rect 178052 388346 178080 404398
rect 181456 402898 181484 405062
rect 183572 405062 184506 405090
rect 181444 402892 181496 402898
rect 181444 402834 181496 402840
rect 179788 399560 179840 399566
rect 179788 399502 179840 399508
rect 178040 388340 178092 388346
rect 178040 388282 178092 388288
rect 178684 388340 178736 388346
rect 178684 388282 178736 388288
rect 178052 387938 178080 388282
rect 178040 387932 178092 387938
rect 178040 387874 178092 387880
rect 178696 381614 178724 388282
rect 178684 381608 178736 381614
rect 178684 381550 178736 381556
rect 177946 380352 178002 380361
rect 177946 380287 178002 380296
rect 177960 310049 177988 380287
rect 178684 369164 178736 369170
rect 178684 369106 178736 369112
rect 178696 363662 178724 369106
rect 179236 364404 179288 364410
rect 179236 364346 179288 364352
rect 178684 363656 178736 363662
rect 178684 363598 178736 363604
rect 178776 357604 178828 357610
rect 178776 357546 178828 357552
rect 178684 357536 178736 357542
rect 178684 357478 178736 357484
rect 177946 310040 178002 310049
rect 177946 309975 178002 309984
rect 177946 308000 178002 308009
rect 177946 307935 178002 307944
rect 177854 305960 177910 305969
rect 177854 305895 177910 305904
rect 177868 305658 177896 305895
rect 177856 305652 177908 305658
rect 177856 305594 177908 305600
rect 177854 301200 177910 301209
rect 177854 301135 177910 301144
rect 177762 270600 177818 270609
rect 177762 270535 177818 270544
rect 177672 225684 177724 225690
rect 177672 225626 177724 225632
rect 177776 160750 177804 270535
rect 177764 160744 177816 160750
rect 177764 160686 177816 160692
rect 177868 151094 177896 301135
rect 177856 151088 177908 151094
rect 177856 151030 177908 151036
rect 177304 146940 177356 146946
rect 177304 146882 177356 146888
rect 177316 110430 177344 146882
rect 177488 118788 177540 118794
rect 177488 118730 177540 118736
rect 177396 113280 177448 113286
rect 177396 113222 177448 113228
rect 177304 110424 177356 110430
rect 177304 110366 177356 110372
rect 177304 103556 177356 103562
rect 177304 103498 177356 103504
rect 177316 90982 177344 103498
rect 177304 90976 177356 90982
rect 177304 90918 177356 90924
rect 177408 86766 177436 113222
rect 177500 93906 177528 118730
rect 177488 93900 177540 93906
rect 177488 93842 177540 93848
rect 177396 86760 177448 86766
rect 177396 86702 177448 86708
rect 176568 25628 176620 25634
rect 176568 25570 176620 25576
rect 175188 20052 175240 20058
rect 175188 19994 175240 20000
rect 177960 10402 177988 307935
rect 178696 257378 178724 357478
rect 178788 352646 178816 357546
rect 178776 352640 178828 352646
rect 178776 352582 178828 352588
rect 179248 341562 179276 364346
rect 179328 363656 179380 363662
rect 179328 363598 179380 363604
rect 179236 341556 179288 341562
rect 179236 341498 179288 341504
rect 179234 292360 179290 292369
rect 179234 292295 179290 292304
rect 179142 263800 179198 263809
rect 179142 263735 179198 263744
rect 178684 257372 178736 257378
rect 178684 257314 178736 257320
rect 178774 256728 178830 256737
rect 178774 256663 178830 256672
rect 178788 226409 178816 256663
rect 178774 226400 178830 226409
rect 178774 226335 178830 226344
rect 178684 109132 178736 109138
rect 178684 109074 178736 109080
rect 178696 79830 178724 109074
rect 179156 91798 179184 263735
rect 179144 91792 179196 91798
rect 179144 91734 179196 91740
rect 179248 84862 179276 292295
rect 179340 286249 179368 363598
rect 179800 352714 179828 399502
rect 181456 394058 181484 402834
rect 181444 394052 181496 394058
rect 181444 393994 181496 394000
rect 183572 373318 183600 405062
rect 187712 399634 187740 405076
rect 187700 399628 187752 399634
rect 187700 399570 187752 399576
rect 190932 396914 190960 405076
rect 193864 402348 193916 402354
rect 193864 402290 193916 402296
rect 190920 396908 190972 396914
rect 190920 396850 190972 396856
rect 183560 373312 183612 373318
rect 183560 373254 183612 373260
rect 190458 365800 190514 365809
rect 190458 365735 190514 365744
rect 190472 364334 190500 365735
rect 190472 364306 191236 364334
rect 187424 360392 187476 360398
rect 187424 360334 187476 360340
rect 181628 358828 181680 358834
rect 181628 358770 181680 358776
rect 181640 355042 181668 358770
rect 182916 357740 182968 357746
rect 182916 357682 182968 357688
rect 181332 355014 181668 355042
rect 182928 355042 182956 357682
rect 184940 357672 184992 357678
rect 184940 357614 184992 357620
rect 184952 355042 184980 357614
rect 187436 355042 187464 360334
rect 189998 360224 190054 360233
rect 189998 360159 190054 360168
rect 190012 355042 190040 360159
rect 182928 355014 183264 355042
rect 184952 355014 185196 355042
rect 187128 355014 187464 355042
rect 189704 355014 190040 355042
rect 191208 355042 191236 364306
rect 193876 359514 193904 402290
rect 194152 398206 194180 405076
rect 197372 404462 197400 405076
rect 200606 405062 200804 405090
rect 197360 404456 197412 404462
rect 197360 404398 197412 404404
rect 197372 402286 197400 404398
rect 200776 402966 200804 405062
rect 203812 404530 203840 405076
rect 202880 404524 202932 404530
rect 202880 404466 202932 404472
rect 203800 404524 203852 404530
rect 203800 404466 203852 404472
rect 200764 402960 200816 402966
rect 200764 402902 200816 402908
rect 197360 402280 197412 402286
rect 197360 402222 197412 402228
rect 194140 398200 194192 398206
rect 194140 398142 194192 398148
rect 194600 398200 194652 398206
rect 194600 398142 194652 398148
rect 193864 359508 193916 359514
rect 193864 359450 193916 359456
rect 193220 356788 193272 356794
rect 193220 356730 193272 356736
rect 193232 355042 193260 356730
rect 194612 355298 194640 398142
rect 200776 370666 200804 402902
rect 202144 395480 202196 395486
rect 202144 395422 202196 395428
rect 200764 370660 200816 370666
rect 200764 370602 200816 370608
rect 197728 359032 197780 359038
rect 197728 358974 197780 358980
rect 194600 355292 194652 355298
rect 194600 355234 194652 355240
rect 195474 355292 195526 355298
rect 195474 355234 195526 355240
rect 191208 355014 191636 355042
rect 193232 355014 193568 355042
rect 179880 354952 179932 354958
rect 179880 354894 179932 354900
rect 179788 352708 179840 352714
rect 179788 352650 179840 352656
rect 179418 343360 179474 343369
rect 179418 343295 179474 343304
rect 179326 286240 179382 286249
rect 179326 286175 179382 286184
rect 179326 268560 179382 268569
rect 179326 268495 179382 268504
rect 179236 84856 179288 84862
rect 179236 84798 179288 84804
rect 178684 79824 178736 79830
rect 178684 79766 178736 79772
rect 179340 26994 179368 268495
rect 179432 243681 179460 343295
rect 179512 341556 179564 341562
rect 179512 341498 179564 341504
rect 179524 341397 179552 341498
rect 179510 341388 179566 341397
rect 179510 341323 179566 341332
rect 179892 274650 179920 354894
rect 194612 354822 194640 355234
rect 195486 355028 195514 355234
rect 197740 355042 197768 358974
rect 202156 358902 202184 395422
rect 202892 365022 202920 404466
rect 206388 399566 206416 405076
rect 209608 402966 209636 405076
rect 212552 405062 212842 405090
rect 215312 405062 216062 405090
rect 218072 405062 219282 405090
rect 222502 405062 222884 405090
rect 209596 402960 209648 402966
rect 209596 402902 209648 402908
rect 206376 399560 206428 399566
rect 206376 399502 206428 399508
rect 212552 392018 212580 405062
rect 214564 401056 214616 401062
rect 214564 400998 214616 401004
rect 212540 392012 212592 392018
rect 212540 391954 212592 391960
rect 212552 391338 212580 391954
rect 212540 391332 212592 391338
rect 212540 391274 212592 391280
rect 205640 373380 205692 373386
rect 205640 373322 205692 373328
rect 202972 371272 203024 371278
rect 202972 371214 203024 371220
rect 202880 365016 202932 365022
rect 202880 364958 202932 364964
rect 202984 364334 203012 371214
rect 205652 367130 205680 373322
rect 209044 371952 209096 371958
rect 209044 371894 209096 371900
rect 205640 367124 205692 367130
rect 205640 367066 205692 367072
rect 205652 364334 205680 367066
rect 209056 364334 209084 371894
rect 211804 367872 211856 367878
rect 211804 367814 211856 367820
rect 202984 364306 203472 364334
rect 205652 364306 206048 364334
rect 202144 358896 202196 358902
rect 202144 358838 202196 358844
rect 199660 356312 199712 356318
rect 199660 356254 199712 356260
rect 199672 355042 199700 356254
rect 202156 355042 202184 358838
rect 197740 355014 198076 355042
rect 199672 355014 200008 355042
rect 201940 355014 202184 355042
rect 203444 355042 203472 364306
rect 206020 355042 206048 364306
rect 208780 364306 209084 364334
rect 208780 357649 208808 364306
rect 208766 357640 208822 357649
rect 211816 357610 211844 367814
rect 208766 357575 208822 357584
rect 211804 357604 211856 357610
rect 208780 355042 208808 357575
rect 211804 357546 211856 357552
rect 211816 355042 211844 357546
rect 214576 356182 214604 400998
rect 215312 371890 215340 405062
rect 217324 378820 217376 378826
rect 217324 378762 217376 378768
rect 217336 371958 217364 378762
rect 218072 378185 218100 405062
rect 222856 404190 222884 405062
rect 224972 405062 225722 405090
rect 227732 405062 228942 405090
rect 222844 404184 222896 404190
rect 222844 404126 222896 404132
rect 218058 378176 218114 378185
rect 218058 378111 218060 378120
rect 218112 378111 218114 378120
rect 218060 378082 218112 378088
rect 220084 376100 220136 376106
rect 220084 376042 220136 376048
rect 217324 371952 217376 371958
rect 217324 371894 217376 371900
rect 215300 371884 215352 371890
rect 215300 371826 215352 371832
rect 220096 358970 220124 376042
rect 220084 358964 220136 358970
rect 220084 358906 220136 358912
rect 220268 358964 220320 358970
rect 220268 358906 220320 358912
rect 217046 358864 217102 358873
rect 217046 358799 217102 358808
rect 214564 356176 214616 356182
rect 214564 356118 214616 356124
rect 214576 355042 214604 356118
rect 217060 355042 217088 358799
rect 218336 357536 218388 357542
rect 218336 357478 218388 357484
rect 203444 355014 203872 355042
rect 206020 355014 206448 355042
rect 208380 355014 208808 355042
rect 209976 355026 210312 355042
rect 209964 355020 210312 355026
rect 210016 355014 210312 355020
rect 211816 355014 212244 355042
rect 214576 355014 214820 355042
rect 216752 355014 217088 355042
rect 218348 355042 218376 357478
rect 220280 355042 220308 358906
rect 222856 355337 222884 404126
rect 224972 393990 225000 405062
rect 224960 393984 225012 393990
rect 224960 393926 225012 393932
rect 227732 370530 227760 405062
rect 232148 402286 232176 405076
rect 234632 405062 235382 405090
rect 236644 405078 236696 405084
rect 232136 402280 232188 402286
rect 232136 402222 232188 402228
rect 234632 385694 234660 405062
rect 234620 385688 234672 385694
rect 234620 385630 234672 385636
rect 234620 383716 234672 383722
rect 234620 383658 234672 383664
rect 231124 373312 231176 373318
rect 231124 373254 231176 373260
rect 227720 370524 227772 370530
rect 227720 370466 227772 370472
rect 225420 358896 225472 358902
rect 225420 358838 225472 358844
rect 223488 357604 223540 357610
rect 223488 357546 223540 357552
rect 222842 355328 222898 355337
rect 222842 355263 222898 355272
rect 223500 355042 223528 357546
rect 225432 355042 225460 358838
rect 227352 357536 227404 357542
rect 227352 357478 227404 357484
rect 227364 355042 227392 357478
rect 228822 356280 228878 356289
rect 228822 356215 228878 356224
rect 218348 355014 218684 355042
rect 220280 355014 220616 355042
rect 223192 355014 223528 355042
rect 225124 355014 225460 355042
rect 227056 355014 227392 355042
rect 209964 354962 210016 354968
rect 194600 354816 194652 354822
rect 194600 354758 194652 354764
rect 228836 354770 228864 356215
rect 231136 356182 231164 373254
rect 234632 364334 234660 383658
rect 236656 376038 236684 405078
rect 237392 405062 238602 405090
rect 241822 405062 242204 405090
rect 236644 376032 236696 376038
rect 236644 375974 236696 375980
rect 237392 369170 237420 405062
rect 242176 404258 242204 405062
rect 242164 404252 242216 404258
rect 242164 404194 242216 404200
rect 239404 403708 239456 403714
rect 239404 403650 239456 403656
rect 239416 370598 239444 403650
rect 240140 403572 240192 403578
rect 240140 403514 240192 403520
rect 240152 396846 240180 403514
rect 240140 396840 240192 396846
rect 240140 396782 240192 396788
rect 241520 394052 241572 394058
rect 241520 393994 241572 394000
rect 239404 370592 239456 370598
rect 239404 370534 239456 370540
rect 237380 369164 237432 369170
rect 237380 369106 237432 369112
rect 234632 364306 235028 364334
rect 233790 359000 233846 359009
rect 233790 358935 233846 358944
rect 231124 356176 231176 356182
rect 231124 356118 231176 356124
rect 231136 355042 231164 356118
rect 233804 355042 233832 358935
rect 231136 355014 231564 355042
rect 233496 355014 233832 355042
rect 235000 355042 235028 364306
rect 237472 362976 237524 362982
rect 237472 362918 237524 362924
rect 240048 362976 240100 362982
rect 240048 362918 240100 362924
rect 235000 355014 235428 355042
rect 237484 354906 237512 362918
rect 240060 355042 240088 362918
rect 239936 355014 240088 355042
rect 241532 355042 241560 393994
rect 242176 384402 242204 404194
rect 242164 384396 242216 384402
rect 242164 384338 242216 384344
rect 242820 363730 242848 405447
rect 242808 363724 242860 363730
rect 242808 363666 242860 363672
rect 242912 360874 242940 532766
rect 242992 532714 243044 532720
rect 243096 532522 243124 538186
rect 243268 532772 243320 532778
rect 243268 532714 243320 532720
rect 243280 532681 243308 532714
rect 243266 532672 243322 532681
rect 243266 532607 243322 532616
rect 243004 532494 243124 532522
rect 243004 400994 243032 532494
rect 243556 407289 243584 580887
rect 244292 409193 244320 700266
rect 244372 630692 244424 630698
rect 244372 630634 244424 630640
rect 244278 409184 244334 409193
rect 244278 409119 244334 409128
rect 243542 407280 243598 407289
rect 243542 407215 243598 407224
rect 243084 407176 243136 407182
rect 243084 407118 243136 407124
rect 243096 405074 243124 407118
rect 243084 405068 243136 405074
rect 243084 405010 243136 405016
rect 242992 400988 243044 400994
rect 242992 400930 243044 400936
rect 243360 369232 243412 369238
rect 243360 369174 243412 369180
rect 243372 368558 243400 369174
rect 242992 368552 243044 368558
rect 242992 368494 243044 368500
rect 243360 368552 243412 368558
rect 243360 368494 243412 368500
rect 243004 364334 243032 368494
rect 243004 364306 243400 364334
rect 242900 360868 242952 360874
rect 242900 360810 242952 360816
rect 243372 355042 243400 364306
rect 244384 359417 244412 630634
rect 245752 599616 245804 599622
rect 245752 599558 245804 599564
rect 244556 594108 244608 594114
rect 244556 594050 244608 594056
rect 244464 588056 244516 588062
rect 244464 587998 244516 588004
rect 244476 403578 244504 587998
rect 244568 515953 244596 594050
rect 245660 585200 245712 585206
rect 245660 585142 245712 585148
rect 245672 583386 245700 585142
rect 245580 583358 245700 583386
rect 245580 582298 245608 583358
rect 245658 583264 245714 583273
rect 245658 583199 245714 583208
rect 245672 582418 245700 583199
rect 245660 582412 245712 582418
rect 245660 582354 245712 582360
rect 245580 582270 245700 582298
rect 244554 515944 244610 515953
rect 244554 515879 244610 515888
rect 245382 515944 245438 515953
rect 245382 515879 245438 515888
rect 245396 514826 245424 515879
rect 245384 514820 245436 514826
rect 245384 514762 245436 514768
rect 245384 447092 245436 447098
rect 245384 447034 245436 447040
rect 245396 445913 245424 447034
rect 244554 445904 244610 445913
rect 244554 445839 244610 445848
rect 245382 445904 245438 445913
rect 245382 445839 245438 445848
rect 244464 403572 244516 403578
rect 244464 403514 244516 403520
rect 244568 367878 244596 445839
rect 245290 409184 245346 409193
rect 245290 409119 245346 409128
rect 245304 408542 245332 409119
rect 245292 408536 245344 408542
rect 245292 408478 245344 408484
rect 245672 407182 245700 582270
rect 245764 576570 245792 599558
rect 245844 595468 245896 595474
rect 245844 595410 245896 595416
rect 245752 576564 245804 576570
rect 245752 576506 245804 576512
rect 245750 576464 245806 576473
rect 245750 576399 245806 576408
rect 245764 575550 245792 576399
rect 245752 575544 245804 575550
rect 245752 575486 245804 575492
rect 245750 573064 245806 573073
rect 245750 572999 245806 573008
rect 245764 572762 245792 572999
rect 245752 572756 245804 572762
rect 245752 572698 245804 572704
rect 245750 566264 245806 566273
rect 245750 566199 245806 566208
rect 245764 565894 245792 566199
rect 245752 565888 245804 565894
rect 245752 565830 245804 565836
rect 245750 560144 245806 560153
rect 245750 560079 245806 560088
rect 245764 558958 245792 560079
rect 245752 558952 245804 558958
rect 245752 558894 245804 558900
rect 245750 556744 245806 556753
rect 245750 556679 245806 556688
rect 245764 556238 245792 556679
rect 245752 556232 245804 556238
rect 245752 556174 245804 556180
rect 245750 549944 245806 549953
rect 245750 549879 245806 549888
rect 245764 549302 245792 549879
rect 245752 549296 245804 549302
rect 245752 549238 245804 549244
rect 245750 539744 245806 539753
rect 245750 539679 245806 539688
rect 245764 539646 245792 539679
rect 245752 539640 245804 539646
rect 245752 539582 245804 539588
rect 245752 539504 245804 539510
rect 245752 539446 245804 539452
rect 245660 407176 245712 407182
rect 245660 407118 245712 407124
rect 245764 384334 245792 539446
rect 245856 536353 245884 595410
rect 246304 587920 246356 587926
rect 246304 587862 246356 587868
rect 245936 576564 245988 576570
rect 245936 576506 245988 576512
rect 245948 569673 245976 576506
rect 245934 569664 245990 569673
rect 245934 569599 245990 569608
rect 245934 543144 245990 543153
rect 245934 543079 245990 543088
rect 245948 539510 245976 543079
rect 245936 539504 245988 539510
rect 245936 539446 245988 539452
rect 245842 536344 245898 536353
rect 245842 536279 245898 536288
rect 245856 536110 245884 536279
rect 245844 536104 245896 536110
rect 245844 536046 245896 536052
rect 245842 526144 245898 526153
rect 245842 526079 245898 526088
rect 245856 525842 245884 526079
rect 245844 525836 245896 525842
rect 245844 525778 245896 525784
rect 245842 522744 245898 522753
rect 245842 522679 245898 522688
rect 245856 521694 245884 522679
rect 245844 521688 245896 521694
rect 245844 521630 245896 521636
rect 245842 519344 245898 519353
rect 245842 519279 245898 519288
rect 245856 518974 245884 519279
rect 245844 518968 245896 518974
rect 245844 518910 245896 518916
rect 245844 512644 245896 512650
rect 245844 512586 245896 512592
rect 245856 512553 245884 512586
rect 245842 512544 245898 512553
rect 245842 512479 245898 512488
rect 245844 506456 245896 506462
rect 245842 506424 245844 506433
rect 245896 506424 245898 506433
rect 245842 506359 245898 506368
rect 245842 503024 245898 503033
rect 245842 502959 245898 502968
rect 245856 502382 245884 502959
rect 245844 502376 245896 502382
rect 245844 502318 245896 502324
rect 245842 499624 245898 499633
rect 245842 499559 245844 499568
rect 245896 499559 245898 499568
rect 245844 499530 245896 499536
rect 245844 496800 245896 496806
rect 245844 496742 245896 496748
rect 245856 496233 245884 496742
rect 245842 496224 245898 496233
rect 245842 496159 245898 496168
rect 245842 492824 245898 492833
rect 245842 492759 245898 492768
rect 245856 492726 245884 492759
rect 245844 492720 245896 492726
rect 245844 492662 245896 492668
rect 245842 486024 245898 486033
rect 245842 485959 245898 485968
rect 245856 485858 245884 485959
rect 245844 485852 245896 485858
rect 245844 485794 245896 485800
rect 245934 479224 245990 479233
rect 245934 479159 245990 479168
rect 245842 475824 245898 475833
rect 245842 475759 245898 475768
rect 245856 474774 245884 475759
rect 245844 474768 245896 474774
rect 245844 474710 245896 474716
rect 245842 472424 245898 472433
rect 245842 472359 245898 472368
rect 245856 472054 245884 472359
rect 245844 472048 245896 472054
rect 245844 471990 245896 471996
rect 245948 470594 245976 479159
rect 245856 470566 245976 470594
rect 245856 395350 245884 470566
rect 245934 462224 245990 462233
rect 245934 462159 245990 462168
rect 245948 460970 245976 462159
rect 245936 460964 245988 460970
rect 245936 460906 245988 460912
rect 245934 459504 245990 459513
rect 245934 459439 245990 459448
rect 245948 458862 245976 459439
rect 245936 458856 245988 458862
rect 245936 458798 245988 458804
rect 245934 456104 245990 456113
rect 245934 456039 245990 456048
rect 245948 455462 245976 456039
rect 245936 455456 245988 455462
rect 245936 455398 245988 455404
rect 246316 450566 246344 587862
rect 247132 583772 247184 583778
rect 247132 583714 247184 583720
rect 246946 562864 247002 562873
rect 247002 562822 247080 562850
rect 246946 562799 247002 562808
rect 246672 509856 246724 509862
rect 246670 509824 246672 509833
rect 246724 509824 246726 509833
rect 246670 509759 246726 509768
rect 246304 450560 246356 450566
rect 246304 450502 246356 450508
rect 245934 449304 245990 449313
rect 245934 449239 245990 449248
rect 245948 448594 245976 449239
rect 245936 448588 245988 448594
rect 245936 448530 245988 448536
rect 246302 442504 246358 442513
rect 246302 442439 246358 442448
rect 245934 439104 245990 439113
rect 245934 439039 245990 439048
rect 245948 438938 245976 439039
rect 245936 438932 245988 438938
rect 245936 438874 245988 438880
rect 245934 435704 245990 435713
rect 245934 435639 245990 435648
rect 245948 434790 245976 435639
rect 245936 434784 245988 434790
rect 245936 434726 245988 434732
rect 245936 433288 245988 433294
rect 245936 433230 245988 433236
rect 245948 432313 245976 433230
rect 245934 432304 245990 432313
rect 245934 432239 245990 432248
rect 245934 428904 245990 428913
rect 245934 428839 245990 428848
rect 245948 427854 245976 428839
rect 245936 427848 245988 427854
rect 245936 427790 245988 427796
rect 245934 425504 245990 425513
rect 245934 425439 245990 425448
rect 245948 425134 245976 425439
rect 245936 425128 245988 425134
rect 245936 425070 245988 425076
rect 245934 422104 245990 422113
rect 245934 422039 245990 422048
rect 245948 420986 245976 422039
rect 245936 420980 245988 420986
rect 245936 420922 245988 420928
rect 245934 418704 245990 418713
rect 245934 418639 245990 418648
rect 245948 418266 245976 418639
rect 245936 418260 245988 418266
rect 245936 418202 245988 418208
rect 245934 415304 245990 415313
rect 245934 415239 245990 415248
rect 245948 414050 245976 415239
rect 245936 414044 245988 414050
rect 245936 413986 245988 413992
rect 245934 411904 245990 411913
rect 245934 411839 245990 411848
rect 245948 411330 245976 411839
rect 245936 411324 245988 411330
rect 245936 411266 245988 411272
rect 245844 395344 245896 395350
rect 245844 395286 245896 395292
rect 246316 393378 246344 442439
rect 246394 405784 246450 405793
rect 246394 405719 246450 405728
rect 246304 393372 246356 393378
rect 246304 393314 246356 393320
rect 246316 392698 246344 393314
rect 246304 392692 246356 392698
rect 246304 392634 246356 392640
rect 246408 392018 246436 405719
rect 246396 392012 246448 392018
rect 246396 391954 246448 391960
rect 246408 391270 246436 391954
rect 246396 391264 246448 391270
rect 246396 391206 246448 391212
rect 245752 384328 245804 384334
rect 245752 384270 245804 384276
rect 247052 376106 247080 562822
rect 247144 482633 247172 583714
rect 248340 509862 248368 702646
rect 283852 702434 283880 703520
rect 297364 702772 297416 702778
rect 297364 702714 297416 702720
rect 282932 702406 283880 702434
rect 253204 700324 253256 700330
rect 253204 700266 253256 700272
rect 251088 643136 251140 643142
rect 251088 643078 251140 643084
rect 249800 588192 249852 588198
rect 249800 588134 249852 588140
rect 248420 586764 248472 586770
rect 248420 586706 248472 586712
rect 248328 509856 248380 509862
rect 248328 509798 248380 509804
rect 248340 509318 248368 509798
rect 248328 509312 248380 509318
rect 248328 509254 248380 509260
rect 247130 482624 247186 482633
rect 247130 482559 247186 482568
rect 247040 376100 247092 376106
rect 247040 376042 247092 376048
rect 244556 367872 244608 367878
rect 244556 367814 244608 367820
rect 245844 363792 245896 363798
rect 245844 363734 245896 363740
rect 244370 359408 244426 359417
rect 244370 359343 244426 359352
rect 241532 355014 241868 355042
rect 243372 355014 243800 355042
rect 237360 354878 237512 354906
rect 245856 354770 245884 363734
rect 247144 356250 247172 482559
rect 247222 465624 247278 465633
rect 247222 465559 247278 465568
rect 247236 395486 247264 465559
rect 247316 418260 247368 418266
rect 247316 418202 247368 418208
rect 247328 401062 247356 418202
rect 248432 403714 248460 586706
rect 248512 558952 248564 558958
rect 248512 558894 248564 558900
rect 248420 403708 248472 403714
rect 248420 403650 248472 403656
rect 247316 401056 247368 401062
rect 247316 400998 247368 401004
rect 247224 395480 247276 395486
rect 247224 395422 247276 395428
rect 248524 377466 248552 558894
rect 249064 456816 249116 456822
rect 249064 456758 249116 456764
rect 249076 404462 249104 456758
rect 249156 407788 249208 407794
rect 249156 407730 249208 407736
rect 249064 404456 249116 404462
rect 249064 404398 249116 404404
rect 249168 402830 249196 407730
rect 249156 402824 249208 402830
rect 249156 402766 249208 402772
rect 249812 395418 249840 588134
rect 251100 512650 251128 643078
rect 251180 591320 251232 591326
rect 251180 591262 251232 591268
rect 251088 512644 251140 512650
rect 251088 512586 251140 512592
rect 249892 509312 249944 509318
rect 249892 509254 249944 509260
rect 249904 405006 249932 509254
rect 251088 482316 251140 482322
rect 251088 482258 251140 482264
rect 249984 458856 250036 458862
rect 249984 458798 250036 458804
rect 249892 405000 249944 405006
rect 249892 404942 249944 404948
rect 249996 403753 250024 458798
rect 251100 433362 251128 482258
rect 251088 433356 251140 433362
rect 251088 433298 251140 433304
rect 249982 403744 250038 403753
rect 249982 403679 250038 403688
rect 249800 395412 249852 395418
rect 249800 395354 249852 395360
rect 251192 378146 251220 591262
rect 252560 586900 252612 586906
rect 252560 586842 252612 586848
rect 251916 585404 251968 585410
rect 251916 585346 251968 585352
rect 251272 583840 251324 583846
rect 251272 583782 251324 583788
rect 251284 403646 251312 583782
rect 251824 510672 251876 510678
rect 251824 510614 251876 510620
rect 251364 425128 251416 425134
rect 251364 425070 251416 425076
rect 251272 403640 251324 403646
rect 251272 403582 251324 403588
rect 251376 398138 251404 425070
rect 251836 404530 251864 510614
rect 251928 485790 251956 585346
rect 251916 485784 251968 485790
rect 251916 485726 251968 485732
rect 252468 425740 252520 425746
rect 252468 425682 252520 425688
rect 252480 425134 252508 425682
rect 252468 425128 252520 425134
rect 252468 425070 252520 425076
rect 251824 404524 251876 404530
rect 251824 404466 251876 404472
rect 251364 398132 251416 398138
rect 251364 398074 251416 398080
rect 251180 378140 251232 378146
rect 251180 378082 251232 378088
rect 252468 378140 252520 378146
rect 252468 378082 252520 378088
rect 252480 377466 252508 378082
rect 248512 377460 248564 377466
rect 248512 377402 248564 377408
rect 252468 377460 252520 377466
rect 252468 377402 252520 377408
rect 252572 369238 252600 586842
rect 252652 450560 252704 450566
rect 252652 450502 252704 450508
rect 252664 402354 252692 450502
rect 252652 402348 252704 402354
rect 252652 402290 252704 402296
rect 253216 373386 253244 700266
rect 262128 698964 262180 698970
rect 262128 698906 262180 698912
rect 256608 594108 256660 594114
rect 256608 594050 256660 594056
rect 255320 586696 255372 586702
rect 255320 586638 255372 586644
rect 253938 583808 253994 583817
rect 253938 583743 253994 583752
rect 253952 387025 253980 583743
rect 255332 400926 255360 586638
rect 255412 448588 255464 448594
rect 255412 448530 255464 448536
rect 255320 400920 255372 400926
rect 255320 400862 255372 400868
rect 253938 387016 253994 387025
rect 253938 386951 253994 386960
rect 255424 381546 255452 448530
rect 256620 402966 256648 594050
rect 258080 589348 258132 589354
rect 258080 589290 258132 589296
rect 256700 588600 256752 588606
rect 256700 588542 256752 588548
rect 256712 588130 256740 588542
rect 256700 588124 256752 588130
rect 256700 588066 256752 588072
rect 256608 402960 256660 402966
rect 256608 402902 256660 402908
rect 256620 402354 256648 402902
rect 256608 402348 256660 402354
rect 256608 402290 256660 402296
rect 256712 398206 256740 588066
rect 257344 536852 257396 536858
rect 257344 536794 257396 536800
rect 257356 404190 257384 536794
rect 257344 404184 257396 404190
rect 257344 404126 257396 404132
rect 256700 398200 256752 398206
rect 256700 398142 256752 398148
rect 258092 392630 258120 589290
rect 260838 586664 260894 586673
rect 260838 586599 260894 586608
rect 259460 586560 259512 586566
rect 259460 586502 259512 586508
rect 258080 392624 258132 392630
rect 258080 392566 258132 392572
rect 256700 391332 256752 391338
rect 256700 391274 256752 391280
rect 255412 381540 255464 381546
rect 255412 381482 255464 381488
rect 253204 373380 253256 373386
rect 253204 373322 253256 373328
rect 252560 369232 252612 369238
rect 252560 369174 252612 369180
rect 250536 360460 250588 360466
rect 250536 360402 250588 360408
rect 247132 356244 247184 356250
rect 247132 356186 247184 356192
rect 247960 356244 248012 356250
rect 247960 356186 248012 356192
rect 247972 355042 248000 356186
rect 250548 355042 250576 360402
rect 254214 357640 254270 357649
rect 254214 357575 254270 357584
rect 254228 356726 254256 357575
rect 254216 356720 254268 356726
rect 254216 356662 254268 356668
rect 252466 356416 252522 356425
rect 252466 356351 252522 356360
rect 252480 355042 252508 356351
rect 247972 355014 248308 355042
rect 250240 355014 250576 355042
rect 252172 355014 252508 355042
rect 254228 354906 254256 356662
rect 256712 355314 256740 391274
rect 259472 367169 259500 586502
rect 259552 518968 259604 518974
rect 259552 518910 259604 518916
rect 259564 399498 259592 518910
rect 260852 405142 260880 586599
rect 262140 496874 262168 698906
rect 278044 697604 278096 697610
rect 278044 697546 278096 697552
rect 263692 585268 263744 585274
rect 263692 585210 263744 585216
rect 263600 514820 263652 514826
rect 263600 514762 263652 514768
rect 262128 496868 262180 496874
rect 262128 496810 262180 496816
rect 261484 485852 261536 485858
rect 261484 485794 261536 485800
rect 260840 405136 260892 405142
rect 260840 405078 260892 405084
rect 259552 399492 259604 399498
rect 259552 399434 259604 399440
rect 261496 373318 261524 485794
rect 263612 390017 263640 514762
rect 263704 506462 263732 585210
rect 276020 581664 276072 581670
rect 276020 581606 276072 581612
rect 264980 549908 265032 549914
rect 264980 549850 265032 549856
rect 264992 549302 265020 549850
rect 264980 549296 265032 549302
rect 264980 549238 265032 549244
rect 263692 506456 263744 506462
rect 263692 506398 263744 506404
rect 263704 505782 263732 506398
rect 263692 505776 263744 505782
rect 263692 505718 263744 505724
rect 263692 455456 263744 455462
rect 263692 455398 263744 455404
rect 263598 390008 263654 390017
rect 263598 389943 263654 389952
rect 262220 384396 262272 384402
rect 262220 384338 262272 384344
rect 261484 373312 261536 373318
rect 261484 373254 261536 373260
rect 259458 367160 259514 367169
rect 259458 367095 259514 367104
rect 260102 367160 260158 367169
rect 260102 367095 260158 367104
rect 260116 358766 260144 367095
rect 260104 358760 260156 358766
rect 260104 358702 260156 358708
rect 260748 357672 260800 357678
rect 260748 357614 260800 357620
rect 258908 356244 258960 356250
rect 258908 356186 258960 356192
rect 254104 354878 254256 354906
rect 256666 355286 256740 355314
rect 256666 354906 256694 355286
rect 258920 355042 258948 356186
rect 260760 355042 260788 357614
rect 262232 357474 262260 384338
rect 263704 367810 263732 455398
rect 264992 374678 265020 549238
rect 270500 492720 270552 492726
rect 270500 492662 270552 492668
rect 269764 460964 269816 460970
rect 269764 460906 269816 460912
rect 264980 374672 265032 374678
rect 264980 374614 265032 374620
rect 264980 370660 265032 370666
rect 264980 370602 265032 370608
rect 263692 367804 263744 367810
rect 263692 367746 263744 367752
rect 262220 357468 262272 357474
rect 262220 357410 262272 357416
rect 256976 355020 257028 355026
rect 258612 355014 258948 355042
rect 260544 355014 260788 355042
rect 262232 355042 262260 357410
rect 264992 355314 265020 370602
rect 269776 367713 269804 460906
rect 270512 378826 270540 492662
rect 275284 470620 275336 470626
rect 275284 470562 275336 470568
rect 275296 382294 275324 470562
rect 273904 382288 273956 382294
rect 273904 382230 273956 382236
rect 275284 382288 275336 382294
rect 275284 382230 275336 382236
rect 271328 379500 271380 379506
rect 271328 379442 271380 379448
rect 271340 378826 271368 379442
rect 270500 378820 270552 378826
rect 270500 378762 270552 378768
rect 271328 378820 271380 378826
rect 271328 378762 271380 378768
rect 270500 377460 270552 377466
rect 270500 377402 270552 377408
rect 269762 367704 269818 367713
rect 269762 367639 269818 367648
rect 266636 358760 266688 358766
rect 266636 358702 266688 358708
rect 264992 355286 265066 355314
rect 262232 355014 262476 355042
rect 265038 355028 265066 355286
rect 266648 355042 266676 358702
rect 270512 355042 270540 377402
rect 273916 364334 273944 382230
rect 276032 365838 276060 581606
rect 278056 447098 278084 697546
rect 282932 592686 282960 702406
rect 291844 670744 291896 670750
rect 291844 670686 291896 670692
rect 282920 592680 282972 592686
rect 282920 592622 282972 592628
rect 289084 587988 289136 587994
rect 289084 587930 289136 587936
rect 287704 572756 287756 572762
rect 287704 572698 287756 572704
rect 282184 525836 282236 525842
rect 282184 525778 282236 525784
rect 278044 447092 278096 447098
rect 278044 447034 278096 447040
rect 278044 438932 278096 438938
rect 278044 438874 278096 438880
rect 278056 377466 278084 438874
rect 278044 377460 278096 377466
rect 278044 377402 278096 377408
rect 282196 371890 282224 525778
rect 287060 377460 287112 377466
rect 287060 377402 287112 377408
rect 279424 371884 279476 371890
rect 279424 371826 279476 371832
rect 282184 371884 282236 371890
rect 282184 371826 282236 371832
rect 276020 365832 276072 365838
rect 276020 365774 276072 365780
rect 273824 364306 273944 364334
rect 276032 364334 276060 365774
rect 276032 364306 276888 364334
rect 273824 355042 273852 364306
rect 266648 355014 266984 355042
rect 270512 355014 270848 355042
rect 273424 355014 273852 355042
rect 276860 355042 276888 364306
rect 279436 357474 279464 371826
rect 287072 364334 287100 377402
rect 287072 364306 287192 364334
rect 282092 357740 282144 357746
rect 282092 357682 282144 357688
rect 279424 357468 279476 357474
rect 279424 357410 279476 357416
rect 279436 355042 279464 357410
rect 282104 355042 282132 357682
rect 276860 355014 277288 355042
rect 279068 355014 279464 355042
rect 281796 355014 282132 355042
rect 283380 355088 283432 355094
rect 287164 355042 287192 364306
rect 287716 362370 287744 572698
rect 287704 362364 287756 362370
rect 287704 362306 287756 362312
rect 289096 356726 289124 587930
rect 291856 425746 291884 670686
rect 292580 585336 292632 585342
rect 292580 585278 292632 585284
rect 291936 427848 291988 427854
rect 291936 427790 291988 427796
rect 291844 425740 291896 425746
rect 291844 425682 291896 425688
rect 291292 365764 291344 365770
rect 291292 365706 291344 365712
rect 290464 357808 290516 357814
rect 290464 357750 290516 357756
rect 289084 356720 289136 356726
rect 289084 356662 289136 356668
rect 290476 355042 290504 357750
rect 283432 355036 283728 355042
rect 283380 355030 283728 355036
rect 283392 355014 283728 355030
rect 287164 355014 287592 355042
rect 290168 355014 290504 355042
rect 256976 354962 257028 354968
rect 256988 354906 257016 354962
rect 256666 354892 257016 354906
rect 256680 354878 257016 354892
rect 279068 354890 279096 355014
rect 287164 354958 287192 355014
rect 287152 354952 287204 354958
rect 285660 354890 285996 354906
rect 287152 354894 287204 354900
rect 279056 354884 279108 354890
rect 285660 354884 286008 354890
rect 285660 354878 285956 354884
rect 279056 354826 279108 354832
rect 285956 354826 286008 354832
rect 269028 354816 269080 354822
rect 228836 354742 228988 354770
rect 245732 354742 245884 354770
rect 268916 354764 269028 354770
rect 268916 354758 269080 354764
rect 268916 354742 269068 354758
rect 275356 354754 275692 354770
rect 275356 354748 275704 354754
rect 275356 354742 275652 354748
rect 275652 354690 275704 354696
rect 291304 354657 291332 365706
rect 291948 364334 291976 427790
rect 292592 368937 292620 585278
rect 296720 512644 296772 512650
rect 296720 512586 296772 512592
rect 292764 414044 292816 414050
rect 292764 413986 292816 413992
rect 292578 368928 292634 368937
rect 292578 368863 292634 368872
rect 292592 368529 292620 368863
rect 292578 368520 292634 368529
rect 292578 368455 292634 368464
rect 291948 364306 292436 364334
rect 291750 357504 291806 357513
rect 291750 357439 291806 357448
rect 291290 354648 291346 354657
rect 291764 354634 291792 357439
rect 292408 354657 292436 364306
rect 292776 356017 292804 413986
rect 293960 387864 294012 387870
rect 293960 387806 294012 387812
rect 293040 387116 293092 387122
rect 293040 387058 293092 387064
rect 292762 356008 292818 356017
rect 292762 355943 292818 355952
rect 292394 354648 292450 354657
rect 291764 354606 292344 354634
rect 291290 354583 291346 354592
rect 292316 354550 292344 354606
rect 292394 354583 292450 354592
rect 292304 354544 292356 354550
rect 292304 354486 292356 354492
rect 293052 350169 293080 387058
rect 293222 368928 293278 368937
rect 293222 368863 293278 368872
rect 293130 356008 293186 356017
rect 293130 355943 293186 355952
rect 293144 354793 293172 355943
rect 293130 354784 293186 354793
rect 293130 354719 293186 354728
rect 293038 350160 293094 350169
rect 293038 350095 293094 350104
rect 293038 347032 293094 347041
rect 293038 346967 293094 346976
rect 179880 274644 179932 274650
rect 179880 274586 179932 274592
rect 179510 262168 179566 262177
rect 179510 262103 179566 262112
rect 179418 243672 179474 243681
rect 179418 243607 179474 243616
rect 179524 243545 179552 262103
rect 179602 244148 179658 244157
rect 179602 244083 179658 244092
rect 179510 243536 179566 243545
rect 179510 243471 179566 243480
rect 179420 242208 179472 242214
rect 179420 242150 179472 242156
rect 179432 239902 179460 242150
rect 179420 239896 179472 239902
rect 179420 239838 179472 239844
rect 179616 238754 179644 244083
rect 215298 240680 215354 240689
rect 190012 240650 190348 240666
rect 190000 240644 190348 240650
rect 190052 240638 190348 240644
rect 215354 240638 215464 240666
rect 292028 240644 292080 240650
rect 215298 240615 215354 240624
rect 190000 240586 190052 240592
rect 292028 240586 292080 240592
rect 287702 240136 287758 240145
rect 180030 239850 180058 240108
rect 179432 238726 179644 238754
rect 179984 239822 180058 239850
rect 180812 240094 181976 240122
rect 183908 240094 184244 240122
rect 179328 26988 179380 26994
rect 179328 26930 179380 26936
rect 179432 14618 179460 238726
rect 179786 231840 179842 231849
rect 179786 231775 179842 231784
rect 179800 231606 179828 231775
rect 179788 231600 179840 231606
rect 179788 231542 179840 231548
rect 179984 219434 180012 239822
rect 179524 219406 180012 219434
rect 179420 14612 179472 14618
rect 179420 14554 179472 14560
rect 179524 11898 179552 219406
rect 180812 32570 180840 240094
rect 184216 237425 184244 240094
rect 184952 240094 185840 240122
rect 184202 237416 184258 237425
rect 184202 237351 184258 237360
rect 184204 187740 184256 187746
rect 184204 187682 184256 187688
rect 184216 158710 184244 187682
rect 184204 158704 184256 158710
rect 184204 158646 184256 158652
rect 184204 151836 184256 151842
rect 184204 151778 184256 151784
rect 182824 140820 182876 140826
rect 182824 140762 182876 140768
rect 181444 139460 181496 139466
rect 181444 139402 181496 139408
rect 181456 92410 181484 139402
rect 182836 93294 182864 140762
rect 182916 118856 182968 118862
rect 182916 118798 182968 118804
rect 182824 93288 182876 93294
rect 182824 93230 182876 93236
rect 181444 92404 181496 92410
rect 181444 92346 181496 92352
rect 182928 89554 182956 118798
rect 184216 90710 184244 151778
rect 184480 140072 184532 140078
rect 184480 140014 184532 140020
rect 184388 124296 184440 124302
rect 184388 124238 184440 124244
rect 184296 110492 184348 110498
rect 184296 110434 184348 110440
rect 184204 90704 184256 90710
rect 184204 90646 184256 90652
rect 182916 89548 182968 89554
rect 182916 89490 182968 89496
rect 184308 77246 184336 110434
rect 184400 90914 184428 124238
rect 184492 109002 184520 140014
rect 184480 108996 184532 109002
rect 184480 108938 184532 108944
rect 184388 90908 184440 90914
rect 184388 90850 184440 90856
rect 184296 77240 184348 77246
rect 184296 77182 184348 77188
rect 184952 75274 184980 240094
rect 187758 239850 187786 240108
rect 187712 239822 187786 239850
rect 191944 240094 192280 240122
rect 193232 240094 194212 240122
rect 195992 240094 196144 240122
rect 186964 207936 187016 207942
rect 186964 207878 187016 207884
rect 185584 191412 185636 191418
rect 185584 191354 185636 191360
rect 185596 95198 185624 191354
rect 185676 147688 185728 147694
rect 185676 147630 185728 147636
rect 185584 95192 185636 95198
rect 185584 95134 185636 95140
rect 185688 88058 185716 147630
rect 185768 117428 185820 117434
rect 185768 117370 185820 117376
rect 185676 88052 185728 88058
rect 185676 87994 185728 88000
rect 185584 87644 185636 87650
rect 185584 87586 185636 87592
rect 184940 75268 184992 75274
rect 184940 75210 184992 75216
rect 180800 32564 180852 32570
rect 180800 32506 180852 32512
rect 179512 11892 179564 11898
rect 179512 11834 179564 11840
rect 177948 10396 178000 10402
rect 177948 10338 178000 10344
rect 175096 4888 175148 4894
rect 175096 4830 175148 4836
rect 185596 3534 185624 87586
rect 185780 75818 185808 117370
rect 186976 95130 187004 207878
rect 187056 137284 187108 137290
rect 187056 137226 187108 137232
rect 186964 95124 187016 95130
rect 186964 95066 187016 95072
rect 187068 92274 187096 137226
rect 187148 98116 187200 98122
rect 187148 98058 187200 98064
rect 187056 92268 187108 92274
rect 187056 92210 187108 92216
rect 187160 81122 187188 98058
rect 187148 81116 187200 81122
rect 187148 81058 187200 81064
rect 185768 75812 185820 75818
rect 185768 75754 185820 75760
rect 187712 17474 187740 239822
rect 191944 237114 191972 240094
rect 191932 237108 191984 237114
rect 191932 237050 191984 237056
rect 192484 235408 192536 235414
rect 192484 235350 192536 235356
rect 189724 225684 189776 225690
rect 189724 225626 189776 225632
rect 188344 176928 188396 176934
rect 188344 176870 188396 176876
rect 188356 171018 188384 176870
rect 188344 171012 188396 171018
rect 188344 170954 188396 170960
rect 188344 128376 188396 128382
rect 188344 128318 188396 128324
rect 188356 79966 188384 128318
rect 188436 121508 188488 121514
rect 188436 121450 188488 121456
rect 188448 85338 188476 121450
rect 188528 107704 188580 107710
rect 188528 107646 188580 107652
rect 188436 85332 188488 85338
rect 188436 85274 188488 85280
rect 188540 81258 188568 107646
rect 188528 81252 188580 81258
rect 188528 81194 188580 81200
rect 188344 79960 188396 79966
rect 188344 79902 188396 79908
rect 187700 17468 187752 17474
rect 187700 17410 187752 17416
rect 189736 3534 189764 225626
rect 191104 183048 191156 183054
rect 191104 182990 191156 182996
rect 189816 127084 189868 127090
rect 189816 127026 189868 127032
rect 189828 78606 189856 127026
rect 189908 111852 189960 111858
rect 189908 111794 189960 111800
rect 189920 82822 189948 111794
rect 189908 82816 189960 82822
rect 189908 82758 189960 82764
rect 191116 82142 191144 182990
rect 191104 82136 191156 82142
rect 191104 82078 191156 82084
rect 189816 78600 189868 78606
rect 189816 78542 189868 78548
rect 192496 7750 192524 235350
rect 192576 184544 192628 184550
rect 192576 184486 192628 184492
rect 192588 91866 192616 184486
rect 192668 160812 192720 160818
rect 192668 160754 192720 160760
rect 192680 150414 192708 160754
rect 192668 150408 192720 150414
rect 192668 150350 192720 150356
rect 192668 138032 192720 138038
rect 192668 137974 192720 137980
rect 192576 91860 192628 91866
rect 192576 91802 192628 91808
rect 192680 78470 192708 137974
rect 192760 106412 192812 106418
rect 192760 106354 192812 106360
rect 192772 81326 192800 106354
rect 192760 81320 192812 81326
rect 192760 81262 192812 81268
rect 192668 78464 192720 78470
rect 192668 78406 192720 78412
rect 192484 7744 192536 7750
rect 192484 7686 192536 7692
rect 193232 4962 193260 240094
rect 195992 238474 196020 240094
rect 198706 239850 198734 240108
rect 200132 240094 200652 240122
rect 201512 240094 202584 240122
rect 204516 240094 204944 240122
rect 198706 239822 198780 239850
rect 195980 238468 196032 238474
rect 195980 238410 196032 238416
rect 195980 238128 196032 238134
rect 195980 238070 196032 238076
rect 195992 233034 196020 238070
rect 195980 233028 196032 233034
rect 195980 232970 196032 232976
rect 198188 227180 198240 227186
rect 198188 227122 198240 227128
rect 196716 217456 196768 217462
rect 196716 217398 196768 217404
rect 196624 190052 196676 190058
rect 196624 189994 196676 190000
rect 195244 151904 195296 151910
rect 195244 151846 195296 151852
rect 193864 139528 193916 139534
rect 193864 139470 193916 139476
rect 193876 86698 193904 139470
rect 194048 104916 194100 104922
rect 194048 104858 194100 104864
rect 193956 96688 194008 96694
rect 193956 96630 194008 96636
rect 193864 86692 193916 86698
rect 193864 86634 193916 86640
rect 193968 84182 193996 96630
rect 194060 94897 194088 104858
rect 194046 94888 194102 94897
rect 194046 94823 194102 94832
rect 195256 94110 195284 151846
rect 195244 94104 195296 94110
rect 195244 94046 195296 94052
rect 193956 84176 194008 84182
rect 193956 84118 194008 84124
rect 196636 9042 196664 189994
rect 196728 185842 196756 217398
rect 198096 187264 198148 187270
rect 198096 187206 198148 187212
rect 196716 185836 196768 185842
rect 196716 185778 196768 185784
rect 196716 180192 196768 180198
rect 196716 180134 196768 180140
rect 196728 90982 196756 180134
rect 198004 177336 198056 177342
rect 198004 177278 198056 177284
rect 196808 120148 196860 120154
rect 196808 120090 196860 120096
rect 196716 90976 196768 90982
rect 196716 90918 196768 90924
rect 196820 82686 196848 120090
rect 196808 82680 196860 82686
rect 196808 82622 196860 82628
rect 196624 9036 196676 9042
rect 196624 8978 196676 8984
rect 198016 6254 198044 177278
rect 198108 82278 198136 187206
rect 198200 177342 198228 227122
rect 198188 177336 198240 177342
rect 198188 177278 198240 177284
rect 198096 82272 198148 82278
rect 198096 82214 198148 82220
rect 198752 6322 198780 239822
rect 199384 113824 199436 113830
rect 199384 113766 199436 113772
rect 199396 95062 199424 113766
rect 199384 95056 199436 95062
rect 199384 94998 199436 95004
rect 200132 31210 200160 240094
rect 200764 110560 200816 110566
rect 200764 110502 200816 110508
rect 200776 86902 200804 110502
rect 200764 86896 200816 86902
rect 200764 86838 200816 86844
rect 201512 32502 201540 240094
rect 204916 238542 204944 240094
rect 207078 239850 207106 240108
rect 209024 240094 209360 240122
rect 207032 239822 207106 239850
rect 204904 238536 204956 238542
rect 204904 238478 204956 238484
rect 203524 221536 203576 221542
rect 203524 221478 203576 221484
rect 203536 184550 203564 221478
rect 204168 191412 204220 191418
rect 204168 191354 204220 191360
rect 203524 184544 203576 184550
rect 203524 184486 203576 184492
rect 202144 153264 202196 153270
rect 202144 153206 202196 153212
rect 202156 92206 202184 153206
rect 203524 146328 203576 146334
rect 203524 146270 203576 146276
rect 202144 92200 202196 92206
rect 202144 92142 202196 92148
rect 203536 85270 203564 146270
rect 203616 114640 203668 114646
rect 203616 114582 203668 114588
rect 203628 88262 203656 114582
rect 203616 88256 203668 88262
rect 203616 88198 203668 88204
rect 203524 85264 203576 85270
rect 203524 85206 203576 85212
rect 201500 32496 201552 32502
rect 201500 32438 201552 32444
rect 200120 31204 200172 31210
rect 200120 31146 200172 31152
rect 198740 6316 198792 6322
rect 198740 6258 198792 6264
rect 198004 6248 198056 6254
rect 198004 6190 198056 6196
rect 193220 4956 193272 4962
rect 193220 4898 193272 4904
rect 204180 3670 204208 191354
rect 204916 155242 204944 238478
rect 206282 177304 206338 177313
rect 206282 177239 206338 177248
rect 204904 155236 204956 155242
rect 204904 155178 204956 155184
rect 204996 153332 205048 153338
rect 204996 153274 205048 153280
rect 204904 102808 204956 102814
rect 204904 102750 204956 102756
rect 204916 3738 204944 102750
rect 205008 94042 205036 153274
rect 205088 107772 205140 107778
rect 205088 107714 205140 107720
rect 204996 94036 205048 94042
rect 204996 93978 205048 93984
rect 205100 79898 205128 107714
rect 205088 79892 205140 79898
rect 205088 79834 205140 79840
rect 206296 6390 206324 177239
rect 206376 150476 206428 150482
rect 206376 150418 206428 150424
rect 206388 111790 206416 150418
rect 206376 111784 206428 111790
rect 206376 111726 206428 111732
rect 206468 104984 206520 104990
rect 206468 104926 206520 104932
rect 206376 103624 206428 103630
rect 206376 103566 206428 103572
rect 206388 86970 206416 103566
rect 206480 93702 206508 104926
rect 206468 93696 206520 93702
rect 206468 93638 206520 93644
rect 206376 86964 206428 86970
rect 206376 86906 206428 86912
rect 207032 17406 207060 239822
rect 209332 237454 209360 240094
rect 210620 240094 210956 240122
rect 212888 240094 213224 240122
rect 210620 238134 210648 240094
rect 210608 238128 210660 238134
rect 210608 238070 210660 238076
rect 213196 237454 213224 240094
rect 216692 240094 217396 240122
rect 218072 240094 219328 240122
rect 220832 240094 221260 240122
rect 223836 240094 224080 240122
rect 209320 237448 209372 237454
rect 209320 237390 209372 237396
rect 210424 237448 210476 237454
rect 210424 237390 210476 237396
rect 213184 237448 213236 237454
rect 213184 237390 213236 237396
rect 216036 237448 216088 237454
rect 216036 237390 216088 237396
rect 209044 179444 209096 179450
rect 209044 179386 209096 179392
rect 209056 165510 209084 179386
rect 209044 165504 209096 165510
rect 209044 165446 209096 165452
rect 209044 142180 209096 142186
rect 209044 142122 209096 142128
rect 207664 138100 207716 138106
rect 207664 138042 207716 138048
rect 207676 92478 207704 138042
rect 207756 111920 207808 111926
rect 207756 111862 207808 111868
rect 207664 92472 207716 92478
rect 207664 92414 207716 92420
rect 207768 74526 207796 111862
rect 209056 82754 209084 142122
rect 209228 102196 209280 102202
rect 209228 102138 209280 102144
rect 209136 99476 209188 99482
rect 209136 99418 209188 99424
rect 209148 89690 209176 99418
rect 209240 93770 209268 102138
rect 209228 93764 209280 93770
rect 209228 93706 209280 93712
rect 209136 89684 209188 89690
rect 209136 89626 209188 89632
rect 209044 82748 209096 82754
rect 209044 82690 209096 82696
rect 207756 74520 207808 74526
rect 207756 74462 207808 74468
rect 210436 25702 210464 237390
rect 214564 234048 214616 234054
rect 214564 233990 214616 233996
rect 211804 214804 211856 214810
rect 211804 214746 211856 214752
rect 211816 178770 211844 214746
rect 214576 190126 214604 233990
rect 214564 190120 214616 190126
rect 214564 190062 214616 190068
rect 214656 189100 214708 189106
rect 214656 189042 214708 189048
rect 211988 180872 212040 180878
rect 211988 180814 212040 180820
rect 211804 178764 211856 178770
rect 211804 178706 211856 178712
rect 211896 178288 211948 178294
rect 211896 178230 211948 178236
rect 211908 164218 211936 178230
rect 212000 168298 212028 180814
rect 214104 179512 214156 179518
rect 214104 179454 214156 179460
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175001 213960 175170
rect 214012 175160 214064 175166
rect 214012 175102 214064 175108
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175102
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 214012 173868 214064 173874
rect 214012 173810 214064 173816
rect 213920 173800 213972 173806
rect 213920 173742 213972 173748
rect 213932 173641 213960 173742
rect 213918 173632 213974 173641
rect 213918 173567 213974 173576
rect 214024 172961 214052 173810
rect 214010 172952 214066 172961
rect 214010 172887 214066 172896
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172281 213960 172450
rect 213918 172272 213974 172281
rect 213918 172207 213974 172216
rect 214116 171601 214144 179454
rect 214564 178152 214616 178158
rect 214564 178094 214616 178100
rect 214102 171592 214158 171601
rect 214102 171527 214158 171536
rect 213920 171080 213972 171086
rect 213918 171048 213920 171057
rect 213972 171048 213974 171057
rect 213918 170983 213974 170992
rect 214012 171012 214064 171018
rect 214012 170954 214064 170960
rect 214024 170377 214052 170954
rect 214010 170368 214066 170377
rect 214010 170303 214066 170312
rect 213920 169720 213972 169726
rect 213920 169662 213972 169668
rect 213932 169017 213960 169662
rect 213918 169008 213974 169017
rect 213918 168943 213974 168952
rect 213920 168360 213972 168366
rect 213920 168302 213972 168308
rect 214010 168328 214066 168337
rect 211988 168292 212040 168298
rect 211988 168234 212040 168240
rect 213932 167657 213960 168302
rect 214010 168263 214012 168272
rect 214064 168263 214066 168272
rect 214012 168234 214064 168240
rect 213918 167648 213974 167657
rect 213918 167583 213974 167592
rect 213920 167000 213972 167006
rect 213918 166968 213920 166977
rect 213972 166968 213974 166977
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 214012 166874 214064 166880
rect 213920 166864 213972 166870
rect 213920 166806 213972 166812
rect 213932 165753 213960 166806
rect 214024 166433 214052 166874
rect 214010 166424 214066 166433
rect 214010 166359 214066 166368
rect 213918 165744 213974 165753
rect 213918 165679 213974 165688
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165073 213960 165514
rect 214012 165504 214064 165510
rect 214012 165446 214064 165452
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214024 164393 214052 165446
rect 214010 164384 214066 164393
rect 214010 164319 214066 164328
rect 211896 164212 211948 164218
rect 211896 164154 211948 164160
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163033 213960 164154
rect 213918 163024 213974 163033
rect 213918 162959 213974 162968
rect 213920 160064 213972 160070
rect 213920 160006 213972 160012
rect 213932 159769 213960 160006
rect 214012 159996 214064 160002
rect 214012 159938 214064 159944
rect 213918 159760 213974 159769
rect 213918 159695 213974 159704
rect 214024 159089 214052 159938
rect 214010 159080 214066 159089
rect 214010 159015 214066 159024
rect 213920 158704 213972 158710
rect 213920 158646 213972 158652
rect 213932 157729 213960 158646
rect 213918 157720 213974 157729
rect 213918 157655 213974 157664
rect 214012 157344 214064 157350
rect 214012 157286 214064 157292
rect 213920 157276 213972 157282
rect 213920 157218 213972 157224
rect 213932 157185 213960 157218
rect 213918 157176 213974 157185
rect 213918 157111 213974 157120
rect 214024 156505 214052 157286
rect 214010 156496 214066 156505
rect 214010 156431 214066 156440
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155825 213960 155858
rect 213918 155816 213974 155825
rect 213918 155751 213974 155760
rect 214010 154456 214066 154465
rect 214010 154391 214066 154400
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 213932 153270 213960 153711
rect 214024 153338 214052 154391
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 214010 153096 214066 153105
rect 214010 153031 214066 153040
rect 213918 152552 213974 152561
rect 213918 152487 213974 152496
rect 213932 151910 213960 152487
rect 213920 151904 213972 151910
rect 213920 151846 213972 151852
rect 214024 151842 214052 153031
rect 214012 151836 214064 151842
rect 214012 151778 214064 151784
rect 214102 151192 214158 151201
rect 214102 151127 214158 151136
rect 211804 151088 211856 151094
rect 211804 151030 211856 151036
rect 210608 127628 210660 127634
rect 210608 127570 210660 127576
rect 210516 121576 210568 121582
rect 210516 121518 210568 121524
rect 210528 84046 210556 121518
rect 210620 93770 210648 127570
rect 210608 93764 210660 93770
rect 210608 93706 210660 93712
rect 210516 84040 210568 84046
rect 210516 83982 210568 83988
rect 210424 25696 210476 25702
rect 210424 25638 210476 25644
rect 207020 17400 207072 17406
rect 207020 17342 207072 17348
rect 206284 6384 206336 6390
rect 206284 6326 206336 6332
rect 211816 3806 211844 151030
rect 213918 150512 213974 150521
rect 213918 150447 213920 150456
rect 213972 150447 213974 150456
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 214024 149161 214052 150350
rect 214010 149152 214066 149161
rect 214010 149087 214066 149096
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148481 213960 148990
rect 213918 148472 213974 148481
rect 213918 148407 213974 148416
rect 213918 147928 213974 147937
rect 213918 147863 213974 147872
rect 213932 147694 213960 147863
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 213918 147248 213974 147257
rect 213918 147183 213974 147192
rect 213932 146334 213960 147183
rect 214116 146946 214144 151127
rect 214576 149841 214604 178094
rect 214668 161809 214696 189042
rect 214932 184952 214984 184958
rect 214932 184894 214984 184900
rect 214840 170400 214892 170406
rect 214840 170342 214892 170348
rect 214654 161800 214710 161809
rect 214654 161735 214710 161744
rect 214852 161474 214880 170342
rect 214944 169697 214972 184894
rect 214930 169688 214986 169697
rect 214930 169623 214986 169632
rect 215024 169040 215076 169046
rect 215024 168982 215076 168988
rect 214852 161446 214972 161474
rect 214944 160449 214972 161446
rect 215036 161129 215064 168982
rect 215022 161120 215078 161129
rect 215022 161055 215078 161064
rect 215944 160744 215996 160750
rect 215944 160686 215996 160692
rect 214930 160440 214986 160449
rect 214930 160375 214986 160384
rect 214654 151872 214710 151881
rect 214654 151807 214710 151816
rect 214562 149832 214618 149841
rect 214562 149767 214618 149776
rect 214104 146940 214156 146946
rect 214104 146882 214156 146888
rect 214562 146568 214618 146577
rect 214562 146503 214618 146512
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 213918 145888 213974 145897
rect 213918 145823 213974 145832
rect 211896 145036 211948 145042
rect 211896 144978 211948 144984
rect 211908 81190 211936 144978
rect 213932 144974 213960 145823
rect 214470 145208 214526 145217
rect 214470 145143 214526 145152
rect 214484 145042 214512 145143
rect 214472 145036 214524 145042
rect 214472 144978 214524 144984
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 213918 144528 213974 144537
rect 213918 144463 213974 144472
rect 213932 143614 213960 144463
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 213918 143304 213974 143313
rect 213918 143239 213974 143248
rect 213932 142186 213960 143239
rect 213920 142180 213972 142186
rect 214576 142154 214604 146503
rect 213920 142122 213972 142128
rect 214484 142126 214604 142154
rect 213918 141944 213974 141953
rect 213918 141879 213974 141888
rect 213182 141264 213238 141273
rect 213182 141199 213238 141208
rect 211988 125724 212040 125730
rect 211988 125666 212040 125672
rect 211896 81184 211948 81190
rect 211896 81126 211948 81132
rect 212000 78538 212028 125666
rect 212080 105052 212132 105058
rect 212080 104994 212132 105000
rect 212092 88330 212120 104994
rect 213196 89622 213224 141199
rect 213932 140826 213960 141879
rect 213920 140820 213972 140826
rect 213920 140762 213972 140768
rect 214010 140584 214066 140593
rect 214010 140519 214066 140528
rect 213918 139904 213974 139913
rect 213918 139839 213974 139848
rect 213932 139466 213960 139839
rect 214024 139534 214052 140519
rect 214012 139528 214064 139534
rect 214012 139470 214064 139476
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 214010 139224 214066 139233
rect 214010 139159 214066 139168
rect 213918 138680 213974 138689
rect 213918 138615 213974 138624
rect 213932 138038 213960 138615
rect 214024 138106 214052 139159
rect 214012 138100 214064 138106
rect 214012 138042 214064 138048
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 214102 138000 214158 138009
rect 214102 137935 214158 137944
rect 214116 136678 214144 137935
rect 214484 137290 214512 142126
rect 214668 140078 214696 151807
rect 214930 142624 214986 142633
rect 214930 142559 214986 142568
rect 214656 140072 214708 140078
rect 214656 140014 214708 140020
rect 214654 137320 214710 137329
rect 214472 137284 214524 137290
rect 214654 137255 214710 137264
rect 214472 137226 214524 137232
rect 214104 136672 214156 136678
rect 214010 136640 214066 136649
rect 214104 136614 214156 136620
rect 214010 136575 214066 136584
rect 213918 135960 213974 135969
rect 213918 135895 213974 135904
rect 213932 135318 213960 135895
rect 214024 135386 214052 136575
rect 214012 135380 214064 135386
rect 214012 135322 214064 135328
rect 213920 135312 213972 135318
rect 213920 135254 213972 135260
rect 214562 135280 214618 135289
rect 214562 135215 214618 135224
rect 213918 134600 213974 134609
rect 213918 134535 213974 134544
rect 213932 133958 213960 134535
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 213918 132696 213974 132705
rect 213918 132631 213974 132640
rect 213932 132530 213960 132631
rect 213920 132524 213972 132530
rect 213920 132466 213972 132472
rect 214010 130656 214066 130665
rect 214010 130591 214066 130600
rect 213918 129976 213974 129985
rect 213918 129911 213974 129920
rect 213932 129878 213960 129911
rect 213920 129872 213972 129878
rect 213920 129814 213972 129820
rect 214024 129810 214052 130591
rect 214012 129804 214064 129810
rect 214012 129746 214064 129752
rect 213918 129296 213974 129305
rect 213918 129231 213974 129240
rect 213932 128382 213960 129231
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 214010 128072 214066 128081
rect 214010 128007 214066 128016
rect 213918 127392 213974 127401
rect 213918 127327 213974 127336
rect 213932 127090 213960 127327
rect 213920 127084 213972 127090
rect 213920 127026 213972 127032
rect 214024 127022 214052 128007
rect 214012 127016 214064 127022
rect 214012 126958 214064 126964
rect 213918 126712 213974 126721
rect 213918 126647 213974 126656
rect 213932 125662 213960 126647
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 125352 214066 125361
rect 214010 125287 214066 125296
rect 213918 124672 213974 124681
rect 213918 124607 213974 124616
rect 213932 124234 213960 124607
rect 214024 124302 214052 125287
rect 214012 124296 214064 124302
rect 214012 124238 214064 124244
rect 213920 124228 213972 124234
rect 213920 124170 213972 124176
rect 214010 124128 214066 124137
rect 214010 124063 214066 124072
rect 213918 123448 213974 123457
rect 213918 123383 213974 123392
rect 213932 122874 213960 123383
rect 214024 122942 214052 124063
rect 214012 122936 214064 122942
rect 214012 122878 214064 122884
rect 213920 122868 213972 122874
rect 213920 122810 213972 122816
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121514 213960 122023
rect 214024 121582 214052 122703
rect 214012 121576 214064 121582
rect 214012 121518 214064 121524
rect 213920 121508 213972 121514
rect 213920 121450 213972 121456
rect 213274 121408 213330 121417
rect 213274 121343 213330 121352
rect 213184 89616 213236 89622
rect 213184 89558 213236 89564
rect 212080 88324 212132 88330
rect 212080 88266 212132 88272
rect 213288 86834 213316 121343
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120154 213960 120663
rect 213920 120148 213972 120154
rect 213920 120090 213972 120096
rect 214102 120048 214158 120057
rect 214102 119983 214158 119992
rect 214010 119504 214066 119513
rect 214010 119439 214066 119448
rect 213920 118856 213972 118862
rect 213918 118824 213920 118833
rect 213972 118824 213974 118833
rect 214024 118794 214052 119439
rect 213918 118759 213974 118768
rect 214012 118788 214064 118794
rect 214012 118730 214064 118736
rect 214116 118726 214144 119983
rect 214104 118720 214156 118726
rect 214104 118662 214156 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 214024 117434 214052 118079
rect 213918 117399 213974 117408
rect 214012 117428 214064 117434
rect 213932 117366 213960 117399
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213920 117302 213972 117308
rect 214010 116784 214066 116793
rect 214010 116719 214066 116728
rect 213918 116104 213974 116113
rect 214024 116074 214052 116719
rect 213918 116039 213974 116048
rect 214012 116068 214064 116074
rect 213932 116006 213960 116039
rect 214012 116010 214064 116016
rect 213920 116000 213972 116006
rect 213920 115942 213972 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114578 213960 114815
rect 214024 114646 214052 115359
rect 214012 114640 214064 114646
rect 214012 114582 214064 114588
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 214010 114200 214066 114209
rect 214010 114135 214066 114144
rect 213918 113520 213974 113529
rect 213918 113455 213974 113464
rect 213932 113286 213960 113455
rect 213920 113280 213972 113286
rect 213920 113222 213972 113228
rect 214024 113218 214052 114135
rect 214012 113212 214064 113218
rect 214012 113154 214064 113160
rect 214010 112840 214066 112849
rect 214010 112775 214066 112784
rect 213918 112160 213974 112169
rect 213918 112095 213974 112104
rect 213932 111858 213960 112095
rect 214024 111926 214052 112775
rect 214012 111920 214064 111926
rect 214012 111862 214064 111868
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110498 213960 110735
rect 214024 110566 214052 111415
rect 214012 110560 214064 110566
rect 214012 110502 214064 110508
rect 213920 110492 213972 110498
rect 213920 110434 213972 110440
rect 214010 110256 214066 110265
rect 214010 110191 214066 110200
rect 213918 109576 213974 109585
rect 213918 109511 213974 109520
rect 213932 109070 213960 109511
rect 214024 109138 214052 110191
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107778 213960 108151
rect 213920 107772 213972 107778
rect 213920 107714 213972 107720
rect 214024 107710 214052 108831
rect 214012 107704 214064 107710
rect 214012 107646 214064 107652
rect 214010 107536 214066 107545
rect 214010 107471 214066 107480
rect 213918 106856 213974 106865
rect 213918 106791 213974 106800
rect 213932 106418 213960 106791
rect 213920 106412 213972 106418
rect 213920 106354 213972 106360
rect 214024 106350 214052 107471
rect 214012 106344 214064 106350
rect 214012 106286 214064 106292
rect 214102 106176 214158 106185
rect 214102 106111 214158 106120
rect 214010 105632 214066 105641
rect 214010 105567 214066 105576
rect 213920 104984 213972 104990
rect 213918 104952 213920 104961
rect 213972 104952 213974 104961
rect 214024 104922 214052 105567
rect 214116 105058 214144 106111
rect 214104 105052 214156 105058
rect 214104 104994 214156 105000
rect 213918 104887 213974 104896
rect 214012 104916 214064 104922
rect 214012 104858 214064 104864
rect 214010 104272 214066 104281
rect 214010 104207 214066 104216
rect 214024 103630 214052 104207
rect 214012 103624 214064 103630
rect 213918 103592 213974 103601
rect 214012 103566 214064 103572
rect 213918 103527 213920 103536
rect 213972 103527 213974 103536
rect 214576 103514 214604 135215
rect 213920 103498 213972 103504
rect 214392 103486 214604 103514
rect 213918 102232 213974 102241
rect 213918 102167 213920 102176
rect 213972 102167 213974 102176
rect 213920 102138 213972 102144
rect 213918 101008 213974 101017
rect 213918 100943 213974 100952
rect 213932 100774 213960 100943
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214010 100328 214066 100337
rect 214010 100263 214066 100272
rect 213918 99648 213974 99657
rect 213918 99583 213974 99592
rect 213932 99414 213960 99583
rect 214024 99482 214052 100263
rect 214012 99476 214064 99482
rect 214012 99418 214064 99424
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214010 98968 214066 98977
rect 214010 98903 214066 98912
rect 213918 98288 213974 98297
rect 213918 98223 213974 98232
rect 213932 98122 213960 98223
rect 213920 98116 213972 98122
rect 213920 98058 213972 98064
rect 214024 98054 214052 98903
rect 214012 98048 214064 98054
rect 214012 97990 214064 97996
rect 213918 97608 213974 97617
rect 213918 97543 213974 97552
rect 213932 96694 213960 97543
rect 214392 97209 214420 103486
rect 214668 101454 214696 137255
rect 214838 132016 214894 132025
rect 214838 131951 214894 131960
rect 214746 126032 214802 126041
rect 214746 125967 214802 125976
rect 214760 125730 214788 125967
rect 214748 125724 214800 125730
rect 214748 125666 214800 125672
rect 214852 122834 214880 131951
rect 214760 122806 214880 122834
rect 214760 122126 214788 122806
rect 214748 122120 214800 122126
rect 214748 122062 214800 122068
rect 214944 120766 214972 142559
rect 214932 120760 214984 120766
rect 214932 120702 214984 120708
rect 214746 102912 214802 102921
rect 214746 102847 214802 102856
rect 214656 101448 214708 101454
rect 214656 101390 214708 101396
rect 214378 97200 214434 97209
rect 214378 97135 214434 97144
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 214654 96384 214710 96393
rect 214654 96319 214710 96328
rect 214562 89176 214618 89185
rect 214562 89111 214618 89120
rect 213276 86828 213328 86834
rect 213276 86770 213328 86776
rect 211988 78532 212040 78538
rect 211988 78474 212040 78480
rect 211804 3800 211856 3806
rect 211804 3742 211856 3748
rect 204904 3732 204956 3738
rect 204904 3674 204956 3680
rect 204168 3664 204220 3670
rect 204168 3606 204220 3612
rect 185584 3528 185636 3534
rect 185584 3470 185636 3476
rect 189724 3528 189776 3534
rect 189724 3470 189776 3476
rect 214576 3466 214604 89111
rect 214668 84114 214696 96319
rect 214760 89729 214788 102847
rect 214930 101552 214986 101561
rect 214930 101487 214986 101496
rect 214838 96928 214894 96937
rect 214838 96863 214894 96872
rect 214746 89720 214802 89729
rect 214746 89655 214802 89664
rect 214852 85542 214880 96863
rect 214944 91050 214972 101487
rect 214932 91044 214984 91050
rect 214932 90986 214984 90992
rect 214840 85536 214892 85542
rect 214840 85478 214892 85484
rect 214656 84108 214708 84114
rect 214656 84050 214708 84056
rect 215956 3466 215984 160686
rect 216048 82210 216076 237390
rect 216128 155236 216180 155242
rect 216128 155178 216180 155184
rect 216036 82204 216088 82210
rect 216036 82146 216088 82152
rect 216140 20670 216168 155178
rect 216692 35290 216720 240094
rect 218072 227662 218100 240094
rect 218060 227656 218112 227662
rect 218060 227598 218112 227604
rect 220084 218884 220136 218890
rect 220084 218826 220136 218832
rect 220096 177410 220124 218826
rect 220832 191418 220860 240094
rect 224052 238785 224080 240094
rect 224972 240094 225768 240122
rect 224038 238776 224094 238785
rect 224038 238711 224094 238720
rect 222844 231192 222896 231198
rect 222844 231134 222896 231140
rect 222856 196858 222884 231134
rect 224224 212016 224276 212022
rect 224224 211958 224276 211964
rect 222844 196852 222896 196858
rect 222844 196794 222896 196800
rect 220820 191412 220872 191418
rect 220820 191354 220872 191360
rect 224236 183054 224264 211958
rect 224972 191185 225000 240094
rect 227686 239850 227714 240108
rect 229112 240094 229632 240122
rect 231872 240094 232208 240122
rect 233896 240094 234140 240122
rect 227686 239822 227760 239850
rect 227732 192778 227760 239822
rect 227720 192772 227772 192778
rect 227720 192714 227772 192720
rect 224958 191176 225014 191185
rect 224958 191111 225014 191120
rect 229112 188601 229140 240094
rect 231872 227118 231900 240094
rect 233896 237114 233924 240094
rect 236058 239850 236086 240108
rect 236012 239822 236086 239850
rect 237392 240094 238004 240122
rect 240580 240094 240824 240122
rect 233884 237108 233936 237114
rect 233884 237050 233936 237056
rect 233896 230382 233924 237050
rect 236012 231606 236040 239822
rect 236000 231600 236052 231606
rect 236000 231542 236052 231548
rect 233884 230376 233936 230382
rect 233884 230318 233936 230324
rect 232504 227248 232556 227254
rect 232504 227190 232556 227196
rect 231860 227112 231912 227118
rect 231860 227054 231912 227060
rect 231124 193996 231176 194002
rect 231124 193938 231176 193944
rect 229098 188592 229154 188601
rect 229098 188527 229154 188536
rect 224224 183048 224276 183054
rect 224224 182990 224276 182996
rect 231136 178945 231164 193938
rect 232516 181694 232544 227190
rect 235264 216164 235316 216170
rect 235264 216106 235316 216112
rect 233884 209228 233936 209234
rect 233884 209170 233936 209176
rect 232504 181688 232556 181694
rect 232504 181630 232556 181636
rect 231122 178936 231178 178945
rect 231122 178871 231178 178880
rect 233896 177478 233924 209170
rect 233976 207868 234028 207874
rect 233976 207810 234028 207816
rect 233988 180198 234016 207810
rect 233976 180192 234028 180198
rect 233976 180134 234028 180140
rect 233884 177472 233936 177478
rect 233884 177414 233936 177420
rect 220084 177404 220136 177410
rect 220084 177346 220136 177352
rect 235276 176662 235304 216106
rect 237392 190058 237420 240094
rect 240796 238542 240824 240094
rect 241532 240094 242512 240122
rect 244292 240094 244444 240122
rect 245672 240094 246376 240122
rect 248432 240094 248952 240122
rect 250548 240094 250884 240122
rect 252816 240094 253060 240122
rect 240784 238536 240836 238542
rect 240784 238478 240836 238484
rect 239496 236700 239548 236706
rect 239496 236642 239548 236648
rect 239404 224256 239456 224262
rect 239404 224198 239456 224204
rect 237380 190052 237432 190058
rect 237380 189994 237432 190000
rect 239416 178809 239444 224198
rect 239508 219434 239536 236642
rect 240796 230314 240824 238478
rect 240784 230308 240836 230314
rect 240784 230250 240836 230256
rect 241532 228954 241560 240094
rect 241520 228948 241572 228954
rect 241520 228890 241572 228896
rect 240784 225616 240836 225622
rect 240784 225558 240836 225564
rect 239496 219428 239548 219434
rect 239496 219370 239548 219376
rect 239496 195492 239548 195498
rect 239496 195434 239548 195440
rect 239402 178800 239458 178809
rect 239402 178735 239458 178744
rect 239508 177614 239536 195434
rect 240796 181762 240824 225558
rect 242164 203652 242216 203658
rect 242164 203594 242216 203600
rect 240784 181756 240836 181762
rect 240784 181698 240836 181704
rect 242176 180334 242204 203594
rect 242256 199572 242308 199578
rect 242256 199514 242308 199520
rect 242164 180328 242216 180334
rect 242164 180270 242216 180276
rect 242268 178022 242296 199514
rect 242348 191344 242400 191350
rect 242348 191286 242400 191292
rect 242360 178838 242388 191286
rect 244292 180266 244320 240094
rect 244924 235340 244976 235346
rect 244924 235282 244976 235288
rect 244936 180402 244964 235282
rect 245672 207874 245700 240094
rect 247684 235272 247736 235278
rect 247684 235214 247736 235220
rect 245660 207868 245712 207874
rect 245660 207810 245712 207816
rect 246304 207800 246356 207806
rect 246304 207742 246356 207748
rect 244924 180396 244976 180402
rect 244924 180338 244976 180344
rect 244280 180260 244332 180266
rect 244280 180202 244332 180208
rect 242348 178832 242400 178838
rect 242348 178774 242400 178780
rect 242256 178016 242308 178022
rect 242256 177958 242308 177964
rect 239496 177608 239548 177614
rect 239496 177550 239548 177556
rect 235264 176656 235316 176662
rect 235264 176598 235316 176604
rect 246316 175982 246344 207742
rect 246396 199640 246448 199646
rect 246396 199582 246448 199588
rect 246408 177313 246436 199582
rect 246488 195424 246540 195430
rect 246488 195366 246540 195372
rect 246500 177546 246528 195366
rect 246488 177540 246540 177546
rect 246488 177482 246540 177488
rect 246394 177304 246450 177313
rect 246394 177239 246450 177248
rect 247696 176089 247724 235214
rect 248432 206650 248460 240094
rect 250548 238746 250576 240094
rect 253032 238882 253060 240094
rect 254412 240094 254748 240122
rect 256712 240094 257324 240122
rect 258092 240094 259256 240122
rect 253020 238876 253072 238882
rect 253020 238818 253072 238824
rect 250536 238740 250588 238746
rect 250536 238682 250588 238688
rect 250548 235278 250576 238682
rect 254412 238610 254440 240094
rect 254400 238604 254452 238610
rect 254400 238546 254452 238552
rect 250536 235272 250588 235278
rect 250536 235214 250588 235220
rect 255320 228404 255372 228410
rect 255320 228346 255372 228352
rect 252836 220176 252888 220182
rect 252836 220118 252888 220124
rect 251180 220108 251232 220114
rect 251180 220050 251232 220056
rect 250444 214668 250496 214674
rect 250444 214610 250496 214616
rect 248420 206644 248472 206650
rect 248420 206586 248472 206592
rect 249800 203720 249852 203726
rect 249800 203662 249852 203668
rect 248512 199504 248564 199510
rect 248512 199446 248564 199452
rect 248524 177585 248552 199446
rect 249064 196784 249116 196790
rect 249064 196726 249116 196732
rect 248510 177576 248566 177585
rect 248510 177511 248566 177520
rect 248052 176656 248104 176662
rect 248052 176598 248104 176604
rect 247682 176080 247738 176089
rect 247682 176015 247738 176024
rect 246304 175976 246356 175982
rect 246304 175918 246356 175924
rect 248064 175817 248092 176598
rect 248050 175808 248106 175817
rect 248050 175743 248106 175752
rect 249076 169130 249104 196726
rect 249340 178016 249392 178022
rect 249340 177958 249392 177964
rect 249154 175944 249210 175953
rect 249154 175879 249210 175888
rect 249168 174729 249196 175879
rect 249352 175273 249380 177958
rect 249338 175264 249394 175273
rect 249338 175199 249394 175208
rect 249154 174720 249210 174729
rect 249154 174655 249210 174664
rect 249154 169144 249210 169153
rect 249076 169102 249154 169130
rect 249154 169079 249210 169088
rect 249708 166320 249760 166326
rect 249708 166262 249760 166268
rect 241520 93900 241572 93906
rect 241520 93842 241572 93848
rect 228364 91928 228416 91934
rect 228364 91870 228416 91876
rect 216680 35284 216732 35290
rect 216680 35226 216732 35232
rect 216128 20664 216180 20670
rect 216128 20606 216180 20612
rect 228376 3602 228404 91870
rect 232504 91860 232556 91866
rect 232504 91802 232556 91808
rect 232516 9110 232544 91802
rect 238760 84924 238812 84930
rect 238760 84866 238812 84872
rect 238024 35284 238076 35290
rect 238024 35226 238076 35232
rect 232504 9104 232556 9110
rect 232504 9046 232556 9052
rect 228364 3596 228416 3602
rect 228364 3538 228416 3544
rect 214564 3460 214616 3466
rect 214564 3402 214616 3408
rect 215944 3460 215996 3466
rect 215944 3402 215996 3408
rect 238036 2990 238064 35226
rect 238772 16574 238800 84866
rect 241532 16574 241560 93842
rect 245660 91792 245712 91798
rect 245660 91734 245712 91740
rect 245672 16574 245700 91734
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 245672 16546 245976 16574
rect 235816 2984 235868 2990
rect 235816 2926 235868 2932
rect 238024 2984 238076 2990
rect 238024 2926 238076 2932
rect 235828 480 235856 2926
rect 239324 480 239352 16546
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 240520 480 240548 3470
rect 241716 480 241744 16546
rect 245200 3800 245252 3806
rect 245200 3742 245252 3748
rect 242900 3732 242952 3738
rect 242900 3674 242952 3680
rect 242912 480 242940 3674
rect 244096 3596 244148 3602
rect 244096 3538 244148 3544
rect 244108 480 244136 3538
rect 245212 480 245240 3742
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247592 4956 247644 4962
rect 247592 4898 247644 4904
rect 247604 480 247632 4898
rect 248788 3664 248840 3670
rect 248788 3606 248840 3612
rect 248800 480 248828 3606
rect 249720 3058 249748 166262
rect 249812 139505 249840 203662
rect 249984 189916 250036 189922
rect 249984 189858 250036 189864
rect 249892 181620 249944 181626
rect 249892 181562 249944 181568
rect 249904 149841 249932 181562
rect 249996 169561 250024 189858
rect 250456 186425 250484 214610
rect 250442 186416 250498 186425
rect 250442 186351 250498 186360
rect 249982 169552 250038 169561
rect 249982 169487 250038 169496
rect 250812 152720 250864 152726
rect 250812 152662 250864 152668
rect 250536 152652 250588 152658
rect 250536 152594 250588 152600
rect 249890 149832 249946 149841
rect 249890 149767 249946 149776
rect 249798 139496 249854 139505
rect 249798 139431 249854 139440
rect 250444 136672 250496 136678
rect 250548 136649 250576 152594
rect 250720 138712 250772 138718
rect 250720 138654 250772 138660
rect 250628 136740 250680 136746
rect 250628 136682 250680 136688
rect 250444 136614 250496 136620
rect 250534 136640 250590 136649
rect 250456 49094 250484 136614
rect 250534 136575 250590 136584
rect 250536 100768 250588 100774
rect 250536 100710 250588 100716
rect 250444 49088 250496 49094
rect 250444 49030 250496 49036
rect 250548 26926 250576 100710
rect 250640 62898 250668 136682
rect 250732 93906 250760 138654
rect 250824 138009 250852 152662
rect 251192 140865 251220 220050
rect 251272 217388 251324 217394
rect 251272 217330 251324 217336
rect 251284 151814 251312 217330
rect 251364 206440 251416 206446
rect 251364 206382 251416 206388
rect 251376 156369 251404 206382
rect 252652 192636 252704 192642
rect 252652 192578 252704 192584
rect 251456 180124 251508 180130
rect 251456 180066 251508 180072
rect 251468 158817 251496 180066
rect 252560 178696 252612 178702
rect 252560 178638 252612 178644
rect 252468 173868 252520 173874
rect 252468 173810 252520 173816
rect 252480 173777 252508 173810
rect 252466 173768 252522 173777
rect 252466 173703 252522 173712
rect 251732 172848 251784 172854
rect 251730 172816 251732 172825
rect 251784 172816 251786 172825
rect 251730 172751 251786 172760
rect 252468 172440 252520 172446
rect 252466 172408 252468 172417
rect 252520 172408 252522 172417
rect 252376 172372 252428 172378
rect 252466 172343 252522 172352
rect 252376 172314 252428 172320
rect 252388 171465 252416 172314
rect 252572 171873 252600 178638
rect 252558 171864 252614 171873
rect 252558 171799 252614 171808
rect 252374 171456 252430 171465
rect 252374 171391 252430 171400
rect 252664 171134 252692 192578
rect 252744 175976 252796 175982
rect 252744 175918 252796 175924
rect 252572 171106 252692 171134
rect 251548 170808 251600 170814
rect 251548 170750 251600 170756
rect 251560 170513 251588 170750
rect 251546 170504 251602 170513
rect 251546 170439 251602 170448
rect 252284 170332 252336 170338
rect 252284 170274 252336 170280
rect 252296 170105 252324 170274
rect 252282 170096 252338 170105
rect 252282 170031 252338 170040
rect 252192 169652 252244 169658
rect 252192 169594 252244 169600
rect 252204 168609 252232 169594
rect 252190 168600 252246 168609
rect 252190 168535 252246 168544
rect 252468 168360 252520 168366
rect 252468 168302 252520 168308
rect 252480 167657 252508 168302
rect 252466 167648 252522 167657
rect 252466 167583 252522 167592
rect 252284 167476 252336 167482
rect 252284 167418 252336 167424
rect 252296 167249 252324 167418
rect 252282 167240 252338 167249
rect 252282 167175 252338 167184
rect 252284 166864 252336 166870
rect 252284 166806 252336 166812
rect 252296 166705 252324 166806
rect 252282 166696 252338 166705
rect 252282 166631 252338 166640
rect 251916 166456 251968 166462
rect 251916 166398 251968 166404
rect 251928 166297 251956 166398
rect 251914 166288 251970 166297
rect 251914 166223 251970 166232
rect 252284 166116 252336 166122
rect 252284 166058 252336 166064
rect 252296 165753 252324 166058
rect 252282 165744 252338 165753
rect 252282 165679 252338 165688
rect 252468 165572 252520 165578
rect 252468 165514 252520 165520
rect 252480 165345 252508 165514
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 251548 164484 251600 164490
rect 251548 164426 251600 164432
rect 251560 164393 251588 164426
rect 251546 164384 251602 164393
rect 251546 164319 251602 164328
rect 252468 164212 252520 164218
rect 252468 164154 252520 164160
rect 252100 164144 252152 164150
rect 252100 164086 252152 164092
rect 252112 163033 252140 164086
rect 252480 163985 252508 164154
rect 252466 163976 252522 163985
rect 252466 163911 252522 163920
rect 252098 163024 252154 163033
rect 252098 162959 252154 162968
rect 252468 162852 252520 162858
rect 252468 162794 252520 162800
rect 252480 162489 252508 162794
rect 252466 162480 252522 162489
rect 252466 162415 252522 162424
rect 252466 162072 252522 162081
rect 252466 162007 252522 162016
rect 252480 161974 252508 162007
rect 252468 161968 252520 161974
rect 252468 161910 252520 161916
rect 252466 161528 252522 161537
rect 252572 161514 252600 171106
rect 252522 161486 252600 161514
rect 252466 161463 252522 161472
rect 252466 161120 252522 161129
rect 252466 161055 252468 161064
rect 252520 161055 252522 161064
rect 252468 161026 252520 161032
rect 252468 160948 252520 160954
rect 252468 160890 252520 160896
rect 252480 160177 252508 160890
rect 252756 160585 252784 175918
rect 252848 164490 252876 220118
rect 253940 210588 253992 210594
rect 253940 210530 253992 210536
rect 252836 164484 252888 164490
rect 252836 164426 252888 164432
rect 252834 164248 252890 164257
rect 252834 164183 252890 164192
rect 252742 160576 252798 160585
rect 252742 160511 252798 160520
rect 252466 160168 252522 160177
rect 252466 160103 252522 160112
rect 252468 160064 252520 160070
rect 252468 160006 252520 160012
rect 251916 159996 251968 160002
rect 251916 159938 251968 159944
rect 251928 159225 251956 159938
rect 252480 159633 252508 160006
rect 252466 159624 252522 159633
rect 252466 159559 252522 159568
rect 251914 159216 251970 159225
rect 251914 159151 251970 159160
rect 252848 159066 252876 164183
rect 253572 160132 253624 160138
rect 253572 160074 253624 160080
rect 252572 159038 252876 159066
rect 251454 158808 251510 158817
rect 251454 158743 251510 158752
rect 252466 158264 252522 158273
rect 252572 158250 252600 159038
rect 252522 158222 252600 158250
rect 252466 158199 252522 158208
rect 252560 158024 252612 158030
rect 252560 157966 252612 157972
rect 251548 157344 251600 157350
rect 251548 157286 251600 157292
rect 252466 157312 252522 157321
rect 251560 156913 251588 157286
rect 252466 157247 252468 157256
rect 252520 157247 252522 157256
rect 252468 157218 252520 157224
rect 251546 156904 251602 156913
rect 251546 156839 251602 156848
rect 251362 156360 251418 156369
rect 251362 156295 251418 156304
rect 252466 155952 252522 155961
rect 252376 155916 252428 155922
rect 252466 155887 252522 155896
rect 252376 155858 252428 155864
rect 251732 155236 251784 155242
rect 251732 155178 251784 155184
rect 251548 154488 251600 154494
rect 251548 154430 251600 154436
rect 251560 154057 251588 154430
rect 251546 154048 251602 154057
rect 251546 153983 251602 153992
rect 251744 152153 251772 155178
rect 252388 155009 252416 155858
rect 252480 155854 252508 155887
rect 252468 155848 252520 155854
rect 252468 155790 252520 155796
rect 252374 155000 252430 155009
rect 252374 154935 252430 154944
rect 252008 154556 252060 154562
rect 252008 154498 252060 154504
rect 252020 153513 252048 154498
rect 252466 154456 252522 154465
rect 252466 154391 252468 154400
rect 252520 154391 252522 154400
rect 252468 154362 252520 154368
rect 252006 153504 252062 153513
rect 252006 153439 252062 153448
rect 252284 153196 252336 153202
rect 252284 153138 252336 153144
rect 252296 152697 252324 153138
rect 252466 153096 252522 153105
rect 252572 153082 252600 157966
rect 253480 154624 253532 154630
rect 253480 154566 253532 154572
rect 252522 153054 252600 153082
rect 252466 153031 252522 153040
rect 252282 152688 252338 152697
rect 252282 152623 252338 152632
rect 251824 152584 251876 152590
rect 251824 152526 251876 152532
rect 251730 152144 251786 152153
rect 251730 152079 251786 152088
rect 251284 151786 251404 151814
rect 251272 151292 251324 151298
rect 251272 151234 251324 151240
rect 251284 151201 251312 151234
rect 251270 151192 251326 151201
rect 251270 151127 251326 151136
rect 251272 147280 251324 147286
rect 251272 147222 251324 147228
rect 251284 146985 251312 147222
rect 251270 146976 251326 146985
rect 251270 146911 251326 146920
rect 251376 146577 251404 151786
rect 251732 149660 251784 149666
rect 251732 149602 251784 149608
rect 251744 149297 251772 149602
rect 251730 149288 251786 149297
rect 251730 149223 251786 149232
rect 251548 148436 251600 148442
rect 251548 148378 251600 148384
rect 251560 148345 251588 148378
rect 251546 148336 251602 148345
rect 251546 148271 251602 148280
rect 251362 146568 251418 146577
rect 251362 146503 251418 146512
rect 251730 146296 251786 146305
rect 251730 146231 251786 146240
rect 251546 144120 251602 144129
rect 251546 144055 251602 144064
rect 251560 143682 251588 144055
rect 251548 143676 251600 143682
rect 251548 143618 251600 143624
rect 251744 143177 251772 146231
rect 251730 143168 251786 143177
rect 251730 143103 251786 143112
rect 251178 140856 251234 140865
rect 251178 140791 251234 140800
rect 251180 140480 251232 140486
rect 251178 140448 251180 140457
rect 251232 140448 251234 140457
rect 251178 140383 251234 140392
rect 251732 138780 251784 138786
rect 251732 138722 251784 138728
rect 250810 138000 250866 138009
rect 250810 137935 250866 137944
rect 251272 137760 251324 137766
rect 251272 137702 251324 137708
rect 251284 137601 251312 137702
rect 251270 137592 251326 137601
rect 251270 137527 251326 137536
rect 251744 135697 251772 138722
rect 251730 135688 251786 135697
rect 251730 135623 251786 135632
rect 251272 133884 251324 133890
rect 251272 133826 251324 133832
rect 251284 133385 251312 133826
rect 251270 133376 251326 133385
rect 251270 133311 251326 133320
rect 251732 132456 251784 132462
rect 251732 132398 251784 132404
rect 251744 131481 251772 132398
rect 251730 131472 251786 131481
rect 251730 131407 251786 131416
rect 251836 128466 251864 152526
rect 252466 151736 252522 151745
rect 252376 151700 252428 151706
rect 252466 151671 252522 151680
rect 252376 151642 252428 151648
rect 252388 150793 252416 151642
rect 252480 151638 252508 151671
rect 252468 151632 252520 151638
rect 252468 151574 252520 151580
rect 252374 150784 252430 150793
rect 252374 150719 252430 150728
rect 252468 150408 252520 150414
rect 252468 150350 252520 150356
rect 252480 150249 252508 150350
rect 252466 150240 252522 150249
rect 252466 150175 252522 150184
rect 252468 149048 252520 149054
rect 252468 148990 252520 148996
rect 252480 148889 252508 148990
rect 252466 148880 252522 148889
rect 252466 148815 252522 148824
rect 252376 147756 252428 147762
rect 252376 147698 252428 147704
rect 252100 146192 252152 146198
rect 252100 146134 252152 146140
rect 252112 145081 252140 146134
rect 252388 145625 252416 147698
rect 252468 147620 252520 147626
rect 252468 147562 252520 147568
rect 252480 147529 252508 147562
rect 252466 147520 252522 147529
rect 252466 147455 252522 147464
rect 252468 146260 252520 146266
rect 252468 146202 252520 146208
rect 252480 146033 252508 146202
rect 252466 146024 252522 146033
rect 252466 145959 252522 145968
rect 252374 145616 252430 145625
rect 252374 145551 252430 145560
rect 252098 145072 252154 145081
rect 252098 145007 252154 145016
rect 252468 144900 252520 144906
rect 252468 144842 252520 144848
rect 252100 144832 252152 144838
rect 252100 144774 252152 144780
rect 252112 143721 252140 144774
rect 252480 144673 252508 144842
rect 252466 144664 252522 144673
rect 252466 144599 252522 144608
rect 252098 143712 252154 143721
rect 252098 143647 252154 143656
rect 253388 143608 253440 143614
rect 253388 143550 253440 143556
rect 251916 142860 251968 142866
rect 251916 142802 251968 142808
rect 251744 128438 251864 128466
rect 251744 126313 251772 128438
rect 251824 128308 251876 128314
rect 251824 128250 251876 128256
rect 251836 127265 251864 128250
rect 251822 127256 251878 127265
rect 251822 127191 251878 127200
rect 251730 126304 251786 126313
rect 251548 126268 251600 126274
rect 251730 126239 251786 126248
rect 251548 126210 251600 126216
rect 251272 124092 251324 124098
rect 251272 124034 251324 124040
rect 251284 123049 251312 124034
rect 251560 124001 251588 126210
rect 251546 123992 251602 124001
rect 251546 123927 251602 123936
rect 251824 123480 251876 123486
rect 251824 123422 251876 123428
rect 251270 123040 251326 123049
rect 251270 122975 251326 122984
rect 251732 122664 251784 122670
rect 251732 122606 251784 122612
rect 251744 122097 251772 122606
rect 251730 122088 251786 122097
rect 251730 122023 251786 122032
rect 251732 121304 251784 121310
rect 251732 121246 251784 121252
rect 251744 120601 251772 121246
rect 251730 120592 251786 120601
rect 251730 120527 251786 120536
rect 251456 120012 251508 120018
rect 251456 119954 251508 119960
rect 251468 118833 251496 119954
rect 251454 118824 251510 118833
rect 251454 118759 251510 118768
rect 251732 118652 251784 118658
rect 251732 118594 251784 118600
rect 251744 117881 251772 118594
rect 251730 117872 251786 117881
rect 251730 117807 251786 117816
rect 251272 117292 251324 117298
rect 251272 117234 251324 117240
rect 251284 116929 251312 117234
rect 251270 116920 251326 116929
rect 251270 116855 251326 116864
rect 251548 115932 251600 115938
rect 251548 115874 251600 115880
rect 251180 115660 251232 115666
rect 251180 115602 251232 115608
rect 251192 115025 251220 115602
rect 251560 115433 251588 115874
rect 251546 115424 251602 115433
rect 251546 115359 251602 115368
rect 251178 115016 251234 115025
rect 251178 114951 251234 114960
rect 251732 113008 251784 113014
rect 251732 112950 251784 112956
rect 251744 112713 251772 112950
rect 251730 112704 251786 112713
rect 251730 112639 251786 112648
rect 251640 111444 251692 111450
rect 251640 111386 251692 111392
rect 251652 111217 251680 111386
rect 251638 111208 251694 111217
rect 251638 111143 251694 111152
rect 251548 110356 251600 110362
rect 251548 110298 251600 110304
rect 251560 110265 251588 110298
rect 251546 110256 251602 110265
rect 251546 110191 251602 110200
rect 251836 107794 251864 123422
rect 251928 115977 251956 142802
rect 253296 142180 253348 142186
rect 253296 142122 253348 142128
rect 252468 141976 252520 141982
rect 252468 141918 252520 141924
rect 252480 141817 252508 141918
rect 252466 141808 252522 141817
rect 252466 141743 252522 141752
rect 252374 141536 252430 141545
rect 252374 141471 252430 141480
rect 252100 136536 252152 136542
rect 252100 136478 252152 136484
rect 252112 135289 252140 136478
rect 252192 135992 252244 135998
rect 252192 135934 252244 135940
rect 252098 135280 252154 135289
rect 252098 135215 252154 135224
rect 252204 134178 252232 135934
rect 252284 135176 252336 135182
rect 252284 135118 252336 135124
rect 252296 134337 252324 135118
rect 252282 134328 252338 134337
rect 252282 134263 252338 134272
rect 252112 134150 252232 134178
rect 252008 131776 252060 131782
rect 252008 131718 252060 131724
rect 251914 115968 251970 115977
rect 251914 115903 251970 115912
rect 252020 111761 252048 131718
rect 252112 124817 252140 134150
rect 252388 134042 252416 141471
rect 252834 141400 252890 141409
rect 252834 141335 252890 141344
rect 252848 141137 252876 141335
rect 252834 141128 252890 141137
rect 252834 141063 252890 141072
rect 253202 140040 253258 140049
rect 253202 139975 253258 139984
rect 252468 139392 252520 139398
rect 252468 139334 252520 139340
rect 252480 138553 252508 139334
rect 252466 138544 252522 138553
rect 252466 138479 252522 138488
rect 252468 137964 252520 137970
rect 252468 137906 252520 137912
rect 252480 137057 252508 137906
rect 252466 137048 252522 137057
rect 252466 136983 252522 136992
rect 252468 136604 252520 136610
rect 252468 136546 252520 136552
rect 252480 136241 252508 136546
rect 252466 136232 252522 136241
rect 252466 136167 252522 136176
rect 252468 135244 252520 135250
rect 252468 135186 252520 135192
rect 252480 134745 252508 135186
rect 252466 134736 252522 134745
rect 252466 134671 252522 134680
rect 252204 134014 252416 134042
rect 252204 132433 252232 134014
rect 252468 133816 252520 133822
rect 252466 133784 252468 133793
rect 252520 133784 252522 133793
rect 252376 133748 252428 133754
rect 252466 133719 252522 133728
rect 252376 133690 252428 133696
rect 252388 132841 252416 133690
rect 252374 132832 252430 132841
rect 252374 132767 252430 132776
rect 252190 132424 252246 132433
rect 252190 132359 252246 132368
rect 252284 132388 252336 132394
rect 252284 132330 252336 132336
rect 252296 131889 252324 132330
rect 252282 131880 252338 131889
rect 252282 131815 252338 131824
rect 252284 131096 252336 131102
rect 252284 131038 252336 131044
rect 252296 130121 252324 131038
rect 252376 131028 252428 131034
rect 252376 130970 252428 130976
rect 252388 130529 252416 130970
rect 252468 130960 252520 130966
rect 252466 130928 252468 130937
rect 252520 130928 252522 130937
rect 252466 130863 252522 130872
rect 252374 130520 252430 130529
rect 252374 130455 252430 130464
rect 252282 130112 252338 130121
rect 252282 130047 252338 130056
rect 252468 129736 252520 129742
rect 252468 129678 252520 129684
rect 252376 129668 252428 129674
rect 252376 129610 252428 129616
rect 252284 129600 252336 129606
rect 252284 129542 252336 129548
rect 252296 128625 252324 129542
rect 252388 129169 252416 129610
rect 252480 129577 252508 129678
rect 252466 129568 252522 129577
rect 252466 129503 252522 129512
rect 252374 129160 252430 129169
rect 252374 129095 252430 129104
rect 252282 128616 252338 128625
rect 252282 128551 252338 128560
rect 252468 128240 252520 128246
rect 252466 128208 252468 128217
rect 252520 128208 252522 128217
rect 252376 128172 252428 128178
rect 252466 128143 252522 128152
rect 252376 128114 252428 128120
rect 252388 127673 252416 128114
rect 252374 127664 252430 127673
rect 252374 127599 252430 127608
rect 252192 126948 252244 126954
rect 252192 126890 252244 126896
rect 252204 125769 252232 126890
rect 252468 126744 252520 126750
rect 252466 126712 252468 126721
rect 252520 126712 252522 126721
rect 252466 126647 252522 126656
rect 252190 125760 252246 125769
rect 252190 125695 252246 125704
rect 252466 125352 252522 125361
rect 252466 125287 252522 125296
rect 252480 125118 252508 125287
rect 252468 125112 252520 125118
rect 252468 125054 252520 125060
rect 252192 124908 252244 124914
rect 252192 124850 252244 124856
rect 252098 124808 252154 124817
rect 252098 124743 252154 124752
rect 252100 119876 252152 119882
rect 252100 119818 252152 119824
rect 252112 113174 252140 119818
rect 252204 119241 252232 124850
rect 252468 124636 252520 124642
rect 252468 124578 252520 124584
rect 252480 124409 252508 124578
rect 252466 124400 252522 124409
rect 252466 124335 252522 124344
rect 252468 124160 252520 124166
rect 252468 124102 252520 124108
rect 252480 123457 252508 124102
rect 252466 123448 252522 123457
rect 252466 123383 252522 123392
rect 252468 122800 252520 122806
rect 252468 122742 252520 122748
rect 252376 122732 252428 122738
rect 252376 122674 252428 122680
rect 252388 121553 252416 122674
rect 252480 122505 252508 122742
rect 252466 122496 252522 122505
rect 252466 122431 252522 122440
rect 252374 121544 252430 121553
rect 252374 121479 252430 121488
rect 252376 121440 252428 121446
rect 252376 121382 252428 121388
rect 252388 120193 252416 121382
rect 252468 121372 252520 121378
rect 252468 121314 252520 121320
rect 252480 121145 252508 121314
rect 252466 121136 252522 121145
rect 252466 121071 252522 121080
rect 252374 120184 252430 120193
rect 252374 120119 252430 120128
rect 252284 120080 252336 120086
rect 252284 120022 252336 120028
rect 252296 119649 252324 120022
rect 252282 119640 252338 119649
rect 252282 119575 252338 119584
rect 252190 119232 252246 119241
rect 252190 119167 252246 119176
rect 252468 118584 252520 118590
rect 252468 118526 252520 118532
rect 252480 118289 252508 118526
rect 252466 118280 252522 118289
rect 252466 118215 252522 118224
rect 252284 117904 252336 117910
rect 252284 117846 252336 117852
rect 252296 117337 252324 117846
rect 252282 117328 252338 117337
rect 252282 117263 252338 117272
rect 252468 117224 252520 117230
rect 252468 117166 252520 117172
rect 252480 116385 252508 117166
rect 252466 116376 252522 116385
rect 252466 116311 252522 116320
rect 252468 114504 252520 114510
rect 252466 114472 252468 114481
rect 252520 114472 252522 114481
rect 252376 114436 252428 114442
rect 252466 114407 252522 114416
rect 252376 114378 252428 114384
rect 252388 114073 252416 114378
rect 252468 114368 252520 114374
rect 252468 114310 252520 114316
rect 252374 114064 252430 114073
rect 252374 113999 252430 114008
rect 252480 113529 252508 114310
rect 252466 113520 252522 113529
rect 252466 113455 252522 113464
rect 252112 113146 252232 113174
rect 252100 112668 252152 112674
rect 252100 112610 252152 112616
rect 252112 112169 252140 112610
rect 252098 112160 252154 112169
rect 252098 112095 252154 112104
rect 252100 111784 252152 111790
rect 252006 111752 252062 111761
rect 252100 111726 252152 111732
rect 252006 111687 252062 111696
rect 251916 111104 251968 111110
rect 251916 111046 251968 111052
rect 251744 107766 251864 107794
rect 251744 105097 251772 107766
rect 251824 107636 251876 107642
rect 251824 107578 251876 107584
rect 251836 107001 251864 107578
rect 251822 106992 251878 107001
rect 251822 106927 251878 106936
rect 251730 105088 251786 105097
rect 251730 105023 251786 105032
rect 251364 104168 251416 104174
rect 251364 104110 251416 104116
rect 251180 102808 251232 102814
rect 251178 102776 251180 102785
rect 251232 102776 251234 102785
rect 251178 102711 251234 102720
rect 251272 102740 251324 102746
rect 251272 102682 251324 102688
rect 251180 101992 251232 101998
rect 251180 101934 251232 101940
rect 251192 101425 251220 101934
rect 251178 101416 251234 101425
rect 251178 101351 251234 101360
rect 251180 97980 251232 97986
rect 251180 97922 251232 97928
rect 251192 96665 251220 97922
rect 251178 96656 251234 96665
rect 251178 96591 251234 96600
rect 250720 93900 250772 93906
rect 250720 93842 250772 93848
rect 250628 62892 250680 62898
rect 250628 62834 250680 62840
rect 250536 26920 250588 26926
rect 250536 26862 250588 26868
rect 251192 11014 251220 96591
rect 251180 11008 251232 11014
rect 251180 10950 251232 10956
rect 251284 6914 251312 102682
rect 251376 98977 251404 104110
rect 251928 101833 251956 111046
rect 252112 110809 252140 111726
rect 252098 110800 252154 110809
rect 252098 110735 252154 110744
rect 252100 110424 252152 110430
rect 252100 110366 252152 110372
rect 252112 109313 252140 110366
rect 252098 109304 252154 109313
rect 252098 109239 252154 109248
rect 252008 108996 252060 109002
rect 252008 108938 252060 108944
rect 252020 107953 252048 108938
rect 252204 108361 252232 113146
rect 252376 112464 252428 112470
rect 252376 112406 252428 112412
rect 252190 108352 252246 108361
rect 252190 108287 252246 108296
rect 252006 107944 252062 107953
rect 252006 107879 252062 107888
rect 252100 107568 252152 107574
rect 252100 107510 252152 107516
rect 252112 106593 252140 107510
rect 252098 106584 252154 106593
rect 252098 106519 252154 106528
rect 252008 106276 252060 106282
rect 252008 106218 252060 106224
rect 252020 106049 252048 106218
rect 252284 106140 252336 106146
rect 252284 106082 252336 106088
rect 252006 106040 252062 106049
rect 252006 105975 252062 105984
rect 252192 104712 252244 104718
rect 252190 104680 252192 104689
rect 252244 104680 252246 104689
rect 252190 104615 252246 104624
rect 252296 103193 252324 106082
rect 252388 104145 252416 112406
rect 252466 109848 252522 109857
rect 252466 109783 252522 109792
rect 252480 109546 252508 109783
rect 252468 109540 252520 109546
rect 252468 109482 252520 109488
rect 252468 108928 252520 108934
rect 252466 108896 252468 108905
rect 252520 108896 252522 108905
rect 252466 108831 252522 108840
rect 252466 107536 252522 107545
rect 252466 107471 252468 107480
rect 252520 107471 252522 107480
rect 252468 107442 252520 107448
rect 252468 105800 252520 105806
rect 252468 105742 252520 105748
rect 252480 105641 252508 105742
rect 252466 105632 252522 105641
rect 252466 105567 252522 105576
rect 252468 104848 252520 104854
rect 252468 104790 252520 104796
rect 252374 104136 252430 104145
rect 252374 104071 252430 104080
rect 252480 103737 252508 104790
rect 252466 103728 252522 103737
rect 252466 103663 252522 103672
rect 252468 103488 252520 103494
rect 252468 103430 252520 103436
rect 252282 103184 252338 103193
rect 252282 103119 252338 103128
rect 252480 102241 252508 103430
rect 252466 102232 252522 102241
rect 252466 102167 252522 102176
rect 252468 102128 252520 102134
rect 252468 102070 252520 102076
rect 251914 101824 251970 101833
rect 251914 101759 251970 101768
rect 252192 101448 252244 101454
rect 252192 101390 252244 101396
rect 252008 100700 252060 100706
rect 252008 100642 252060 100648
rect 251548 100564 251600 100570
rect 251548 100506 251600 100512
rect 251560 100473 251588 100506
rect 251546 100464 251602 100473
rect 251546 100399 251602 100408
rect 252020 99929 252048 100642
rect 252006 99920 252062 99929
rect 252006 99855 252062 99864
rect 251362 98968 251418 98977
rect 251362 98903 251418 98912
rect 252204 97073 252232 101390
rect 252480 100881 252508 102070
rect 252466 100872 252522 100881
rect 252466 100807 252522 100816
rect 252468 100632 252520 100638
rect 252468 100574 252520 100580
rect 252480 99521 252508 100574
rect 252466 99512 252522 99521
rect 252466 99447 252522 99456
rect 252468 98864 252520 98870
rect 252468 98806 252520 98812
rect 252480 98569 252508 98806
rect 252466 98560 252522 98569
rect 252466 98495 252522 98504
rect 253216 97986 253244 139975
rect 253308 101998 253336 142122
rect 253400 102814 253428 143550
rect 253492 115666 253520 154566
rect 253584 140486 253612 160074
rect 253952 151298 253980 210530
rect 254032 192704 254084 192710
rect 254032 192646 254084 192652
rect 253940 151292 253992 151298
rect 253940 151234 253992 151240
rect 254044 147286 254072 192646
rect 254216 184408 254268 184414
rect 254216 184350 254268 184356
rect 254122 177304 254178 177313
rect 254122 177239 254178 177248
rect 254032 147280 254084 147286
rect 254032 147222 254084 147228
rect 253572 140480 253624 140486
rect 253572 140422 253624 140428
rect 254136 137766 254164 177239
rect 254228 170814 254256 184350
rect 254216 170808 254268 170814
rect 254216 170750 254268 170756
rect 255332 160138 255360 228346
rect 256712 220114 256740 240094
rect 256700 220108 256752 220114
rect 256700 220050 256752 220056
rect 258092 215422 258120 240094
rect 261174 239850 261202 240108
rect 261128 239822 261202 239850
rect 262232 240094 263120 240122
rect 265544 240094 265696 240122
rect 267292 240094 267628 240122
rect 269224 240094 269560 240122
rect 271156 240094 271492 240122
rect 258080 215416 258132 215422
rect 258080 215358 258132 215364
rect 259460 213376 259512 213382
rect 259460 213318 259512 213324
rect 256976 200932 257028 200938
rect 256976 200874 257028 200880
rect 255412 191276 255464 191282
rect 255412 191218 255464 191224
rect 255320 160132 255372 160138
rect 255320 160074 255372 160080
rect 254676 149728 254728 149734
rect 254676 149670 254728 149676
rect 254584 144968 254636 144974
rect 254584 144910 254636 144916
rect 254124 137760 254176 137766
rect 254124 137702 254176 137708
rect 253480 115660 253532 115666
rect 253480 115602 253532 115608
rect 254596 106146 254624 144910
rect 254688 111450 254716 149670
rect 255424 148442 255452 191218
rect 256792 187060 256844 187066
rect 256792 187002 256844 187008
rect 255596 185768 255648 185774
rect 255596 185710 255648 185716
rect 255504 180396 255556 180402
rect 255504 180338 255556 180344
rect 255516 149666 255544 180338
rect 255608 172854 255636 185710
rect 256700 177608 256752 177614
rect 256700 177550 256752 177556
rect 255596 172848 255648 172854
rect 255596 172790 255648 172796
rect 256712 167482 256740 177550
rect 256804 170338 256832 187002
rect 256884 180328 256936 180334
rect 256884 180270 256936 180276
rect 256792 170332 256844 170338
rect 256792 170274 256844 170280
rect 256790 169824 256846 169833
rect 256790 169759 256846 169768
rect 256700 167476 256752 167482
rect 256700 167418 256752 167424
rect 255964 152516 256016 152522
rect 255964 152458 256016 152464
rect 255504 149660 255556 149666
rect 255504 149602 255556 149608
rect 255412 148436 255464 148442
rect 255412 148378 255464 148384
rect 254768 148368 254820 148374
rect 254768 148310 254820 148316
rect 254780 120018 254808 148310
rect 254768 120012 254820 120018
rect 254768 119954 254820 119960
rect 255976 113014 256004 152458
rect 256332 151088 256384 151094
rect 256332 151030 256384 151036
rect 256240 146396 256292 146402
rect 256240 146338 256292 146344
rect 256148 146328 256200 146334
rect 256148 146270 256200 146276
rect 255964 113008 256016 113014
rect 255964 112950 256016 112956
rect 256056 111852 256108 111858
rect 256056 111794 256108 111800
rect 254676 111444 254728 111450
rect 254676 111386 254728 111392
rect 254584 106140 254636 106146
rect 254584 106082 254636 106088
rect 255964 105596 256016 105602
rect 255964 105538 256016 105544
rect 253388 102808 253440 102814
rect 253388 102750 253440 102756
rect 253296 101992 253348 101998
rect 253296 101934 253348 101940
rect 253204 97980 253256 97986
rect 253204 97922 253256 97928
rect 252190 97064 252246 97073
rect 252190 96999 252246 97008
rect 253296 96688 253348 96694
rect 253296 96630 253348 96636
rect 251362 96248 251418 96257
rect 251362 96183 251418 96192
rect 251376 35290 251404 96183
rect 252560 86284 252612 86290
rect 252560 86226 252612 86232
rect 251364 35284 251416 35290
rect 251364 35226 251416 35232
rect 252572 16574 252600 86226
rect 253308 21418 253336 96630
rect 253296 21412 253348 21418
rect 253296 21354 253348 21360
rect 253204 17468 253256 17474
rect 253204 17410 253256 17416
rect 252572 16546 253152 16574
rect 251192 6886 251312 6914
rect 249984 4956 250036 4962
rect 249984 4898 250036 4904
rect 249708 3052 249760 3058
rect 249708 2994 249760 3000
rect 249996 480 250024 4898
rect 251192 480 251220 6886
rect 252376 3528 252428 3534
rect 252376 3470 252428 3476
rect 253124 3482 253152 16546
rect 253216 3670 253244 17410
rect 253204 3664 253256 3670
rect 253204 3606 253256 3612
rect 255976 3602 256004 105538
rect 256068 14550 256096 111794
rect 256160 104718 256188 146270
rect 256252 105806 256280 146338
rect 256344 112674 256372 151030
rect 256804 141982 256832 169759
rect 256896 166122 256924 180270
rect 256884 166116 256936 166122
rect 256884 166058 256936 166064
rect 256988 147762 257016 200874
rect 258172 189984 258224 189990
rect 258172 189926 258224 189932
rect 258080 178764 258132 178770
rect 258080 178706 258132 178712
rect 258092 173874 258120 178706
rect 258080 173868 258132 173874
rect 258080 173810 258132 173816
rect 258080 173732 258132 173738
rect 258080 173674 258132 173680
rect 258092 169658 258120 173674
rect 258080 169652 258132 169658
rect 258080 169594 258132 169600
rect 258184 166870 258212 189926
rect 258264 181688 258316 181694
rect 258264 181630 258316 181636
rect 258172 166864 258224 166870
rect 258172 166806 258224 166812
rect 257528 165640 257580 165646
rect 257528 165582 257580 165588
rect 257436 157412 257488 157418
rect 257436 157354 257488 157360
rect 256976 147756 257028 147762
rect 256976 147698 257028 147704
rect 257344 147688 257396 147694
rect 257344 147630 257396 147636
rect 256792 141976 256844 141982
rect 256792 141918 256844 141924
rect 256700 130416 256752 130422
rect 256700 130358 256752 130364
rect 256332 112668 256384 112674
rect 256332 112610 256384 112616
rect 256240 105800 256292 105806
rect 256240 105742 256292 105748
rect 256148 104712 256200 104718
rect 256148 104654 256200 104660
rect 256148 98048 256200 98054
rect 256148 97990 256200 97996
rect 256160 17270 256188 97990
rect 256148 17264 256200 17270
rect 256148 17206 256200 17212
rect 256056 14544 256108 14550
rect 256056 14486 256108 14492
rect 255964 3596 256016 3602
rect 255964 3538 256016 3544
rect 252388 480 252416 3470
rect 253124 3454 253520 3482
rect 253492 480 253520 3454
rect 254676 3460 254728 3466
rect 254676 3402 254728 3408
rect 254688 480 254716 3402
rect 255872 3052 255924 3058
rect 255872 2994 255924 3000
rect 255884 480 255912 2994
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 130358
rect 257356 107506 257384 147630
rect 257448 117910 257476 157354
rect 257540 126750 257568 165582
rect 258276 161090 258304 181630
rect 258448 178832 258500 178838
rect 258448 178774 258500 178780
rect 258356 177472 258408 177478
rect 258356 177414 258408 177420
rect 258368 173738 258396 177414
rect 258356 173732 258408 173738
rect 258356 173674 258408 173680
rect 258460 161474 258488 178774
rect 258908 167680 258960 167686
rect 258908 167622 258960 167628
rect 258368 161446 258488 161474
rect 258816 161492 258868 161498
rect 258264 161084 258316 161090
rect 258264 161026 258316 161032
rect 258368 152726 258396 161446
rect 258816 161434 258868 161440
rect 258356 152720 258408 152726
rect 258356 152662 258408 152668
rect 258724 150476 258776 150482
rect 258724 150418 258776 150424
rect 257528 126744 257580 126750
rect 257528 126686 257580 126692
rect 257436 117904 257488 117910
rect 257436 117846 257488 117852
rect 258736 109546 258764 150418
rect 258828 122670 258856 161434
rect 258920 132394 258948 167622
rect 259000 159384 259052 159390
rect 259000 159326 259052 159332
rect 258908 132388 258960 132394
rect 258908 132330 258960 132336
rect 259012 125118 259040 159326
rect 259472 143682 259500 213318
rect 259552 191208 259604 191214
rect 259552 191150 259604 191156
rect 259564 166462 259592 191150
rect 259644 185836 259696 185842
rect 259644 185778 259696 185784
rect 259552 166456 259604 166462
rect 259552 166398 259604 166404
rect 259656 161974 259684 185778
rect 259736 184544 259788 184550
rect 259736 184486 259788 184492
rect 259644 161968 259696 161974
rect 259644 161910 259696 161916
rect 259748 160954 259776 184486
rect 260932 183048 260984 183054
rect 260932 182990 260984 182996
rect 260840 180192 260892 180198
rect 260840 180134 260892 180140
rect 260852 172446 260880 180134
rect 260840 172440 260892 172446
rect 260840 172382 260892 172388
rect 260196 164280 260248 164286
rect 260196 164222 260248 164228
rect 259736 160948 259788 160954
rect 259736 160890 259788 160896
rect 260104 160132 260156 160138
rect 260104 160074 260156 160080
rect 259460 143676 259512 143682
rect 259460 143618 259512 143624
rect 259000 125112 259052 125118
rect 259000 125054 259052 125060
rect 258816 122664 258868 122670
rect 258816 122606 258868 122612
rect 260116 121310 260144 160074
rect 260208 124642 260236 164222
rect 260944 158030 260972 182990
rect 261022 173904 261078 173913
rect 261022 173839 261078 173848
rect 260932 158024 260984 158030
rect 260932 157966 260984 157972
rect 261036 152658 261064 173839
rect 261128 163538 261156 239822
rect 262232 222193 262260 240094
rect 265544 238746 265572 240094
rect 265532 238740 265584 238746
rect 265532 238682 265584 238688
rect 265544 234530 265572 238682
rect 267292 237454 267320 240094
rect 265624 237448 265676 237454
rect 265624 237390 265676 237396
rect 267280 237448 267332 237454
rect 267280 237390 267332 237396
rect 265532 234524 265584 234530
rect 265532 234466 265584 234472
rect 264336 233980 264388 233986
rect 264336 233922 264388 233928
rect 262218 222184 262274 222193
rect 262218 222119 262274 222128
rect 262862 222184 262918 222193
rect 262862 222119 262918 222128
rect 262404 196920 262456 196926
rect 262404 196862 262456 196868
rect 262220 181756 262272 181762
rect 262220 181698 262272 181704
rect 261116 163532 261168 163538
rect 261116 163474 261168 163480
rect 261484 160744 261536 160750
rect 261484 160686 261536 160692
rect 261024 152652 261076 152658
rect 261024 152594 261076 152600
rect 260380 149116 260432 149122
rect 260380 149058 260432 149064
rect 260288 125656 260340 125662
rect 260288 125598 260340 125604
rect 260196 124636 260248 124642
rect 260196 124578 260248 124584
rect 260104 121304 260156 121310
rect 260104 121246 260156 121252
rect 260104 119400 260156 119406
rect 260104 119342 260156 119348
rect 258724 109540 258776 109546
rect 258724 109482 258776 109488
rect 257344 107500 257396 107506
rect 257344 107442 257396 107448
rect 260116 98870 260144 119342
rect 260104 98864 260156 98870
rect 260104 98806 260156 98812
rect 260196 98116 260248 98122
rect 260196 98058 260248 98064
rect 258080 95940 258132 95946
rect 258080 95882 258132 95888
rect 258092 16574 258120 95882
rect 260104 82272 260156 82278
rect 260104 82214 260156 82220
rect 258092 16546 258304 16574
rect 258276 480 258304 16546
rect 260116 6458 260144 82214
rect 260208 44946 260236 98058
rect 260300 91934 260328 125598
rect 260392 119882 260420 149058
rect 261496 129606 261524 160686
rect 261576 155984 261628 155990
rect 261576 155926 261628 155932
rect 261484 129600 261536 129606
rect 261484 129542 261536 129548
rect 261484 121508 261536 121514
rect 261484 121450 261536 121456
rect 260380 119876 260432 119882
rect 260380 119818 260432 119824
rect 260288 91928 260340 91934
rect 260288 91870 260340 91876
rect 260196 44940 260248 44946
rect 260196 44882 260248 44888
rect 261496 28354 261524 121450
rect 261588 117230 261616 155926
rect 261668 153264 261720 153270
rect 261668 153206 261720 153212
rect 261576 117224 261628 117230
rect 261576 117166 261628 117172
rect 261680 114374 261708 153206
rect 261760 145580 261812 145586
rect 261760 145522 261812 145528
rect 261772 122738 261800 145522
rect 262232 144838 262260 181698
rect 262312 177404 262364 177410
rect 262312 177346 262364 177352
rect 262324 151706 262352 177346
rect 262416 172378 262444 196862
rect 262876 174554 262904 222119
rect 264244 215416 264296 215422
rect 264244 215358 264296 215364
rect 263692 188488 263744 188494
rect 263692 188430 263744 188436
rect 263600 177336 263652 177342
rect 263600 177278 263652 177284
rect 262864 174548 262916 174554
rect 262864 174490 262916 174496
rect 262404 172372 262456 172378
rect 262404 172314 262456 172320
rect 262956 171148 263008 171154
rect 262956 171090 263008 171096
rect 262312 151700 262364 151706
rect 262312 151642 262364 151648
rect 262220 144832 262272 144838
rect 262220 144774 262272 144780
rect 262864 141432 262916 141438
rect 262864 141374 262916 141380
rect 261760 122732 261812 122738
rect 261760 122674 261812 122680
rect 261668 114368 261720 114374
rect 261668 114310 261720 114316
rect 261576 106344 261628 106350
rect 261576 106286 261628 106292
rect 261588 64258 261616 106286
rect 262876 103494 262904 141374
rect 262968 133754 262996 171090
rect 263048 162172 263100 162178
rect 263048 162114 263100 162120
rect 262956 133748 263008 133754
rect 262956 133690 263008 133696
rect 263060 128178 263088 162114
rect 263612 155854 263640 177278
rect 263704 168366 263732 188430
rect 263692 168360 263744 168366
rect 263692 168302 263744 168308
rect 263600 155848 263652 155854
rect 263600 155790 263652 155796
rect 263140 133204 263192 133210
rect 263140 133146 263192 133152
rect 263048 128172 263100 128178
rect 263048 128114 263100 128120
rect 262956 116000 263008 116006
rect 262956 115942 263008 115948
rect 262864 103488 262916 103494
rect 262864 103430 262916 103436
rect 261668 102196 261720 102202
rect 261668 102138 261720 102144
rect 261680 71126 261708 102138
rect 262864 96756 262916 96762
rect 262864 96698 262916 96704
rect 261668 71120 261720 71126
rect 261668 71062 261720 71068
rect 261576 64252 261628 64258
rect 261576 64194 261628 64200
rect 261576 32564 261628 32570
rect 261576 32506 261628 32512
rect 261484 28348 261536 28354
rect 261484 28290 261536 28296
rect 260656 9036 260708 9042
rect 260656 8978 260708 8984
rect 260104 6452 260156 6458
rect 260104 6394 260156 6400
rect 259460 3596 259512 3602
rect 259460 3538 259512 3544
rect 259472 480 259500 3538
rect 260668 480 260696 8978
rect 261588 4146 261616 32506
rect 262876 24138 262904 96698
rect 262968 50386 262996 115942
rect 263152 107574 263180 133146
rect 263140 107568 263192 107574
rect 263140 107510 263192 107516
rect 262956 50380 263008 50386
rect 262956 50322 263008 50328
rect 262864 24132 262916 24138
rect 262864 24074 262916 24080
rect 262220 20052 262272 20058
rect 262220 19994 262272 20000
rect 262232 16574 262260 19994
rect 262232 16546 262536 16574
rect 261576 4140 261628 4146
rect 261576 4082 261628 4088
rect 261760 3664 261812 3670
rect 261760 3606 261812 3612
rect 261772 480 261800 3606
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264152 3460 264204 3466
rect 264152 3402 264204 3408
rect 264164 480 264192 3402
rect 264256 3262 264284 215358
rect 264348 191214 264376 233922
rect 264980 203856 265032 203862
rect 264980 203798 265032 203804
rect 264336 191208 264388 191214
rect 264336 191150 264388 191156
rect 264336 168428 264388 168434
rect 264336 168370 264388 168376
rect 264348 129674 264376 168370
rect 264992 164150 265020 203798
rect 264980 164144 265032 164150
rect 264980 164086 265032 164092
rect 264428 157480 264480 157486
rect 264428 157422 264480 157428
rect 264336 129668 264388 129674
rect 264336 129610 264388 129616
rect 264336 124432 264388 124438
rect 264336 124374 264388 124380
rect 264348 13122 264376 124374
rect 264440 118590 264468 157422
rect 264888 135924 264940 135930
rect 264888 135866 264940 135872
rect 264428 118584 264480 118590
rect 264428 118526 264480 118532
rect 264336 13116 264388 13122
rect 264336 13058 264388 13064
rect 264900 3738 264928 135866
rect 264980 117972 265032 117978
rect 264980 117914 265032 117920
rect 264888 3732 264940 3738
rect 264888 3674 264940 3680
rect 264244 3256 264296 3262
rect 264244 3198 264296 3204
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 117914
rect 265636 4962 265664 237390
rect 269224 237182 269252 240094
rect 269212 237176 269264 237182
rect 269212 237118 269264 237124
rect 271156 232966 271184 240094
rect 274054 239850 274082 240108
rect 275986 239850 276014 240108
rect 277412 240094 277932 240122
rect 278884 240094 279864 240122
rect 281552 240094 282440 240122
rect 274054 239822 274128 239850
rect 275986 239822 276060 239850
rect 274100 235890 274128 239822
rect 276032 238678 276060 239822
rect 276020 238672 276072 238678
rect 276020 238614 276072 238620
rect 274088 235884 274140 235890
rect 274088 235826 274140 235832
rect 275282 235376 275338 235385
rect 275282 235311 275338 235320
rect 271144 232960 271196 232966
rect 271144 232902 271196 232908
rect 268384 227112 268436 227118
rect 268384 227054 268436 227060
rect 267832 203788 267884 203794
rect 267832 203730 267884 203736
rect 266360 198212 266412 198218
rect 266360 198154 266412 198160
rect 265900 173936 265952 173942
rect 265900 173878 265952 173884
rect 265716 172576 265768 172582
rect 265716 172518 265768 172524
rect 265728 133822 265756 172518
rect 265808 158772 265860 158778
rect 265808 158714 265860 158720
rect 265716 133816 265768 133822
rect 265716 133758 265768 133764
rect 265716 124296 265768 124302
rect 265716 124238 265768 124244
rect 265728 11830 265756 124238
rect 265820 120086 265848 158714
rect 265912 136542 265940 173878
rect 266372 144906 266400 198154
rect 266452 193928 266504 193934
rect 266452 193870 266504 193876
rect 266464 160002 266492 193870
rect 267740 187196 267792 187202
rect 267740 187138 267792 187144
rect 267188 169788 267240 169794
rect 267188 169730 267240 169736
rect 267096 167068 267148 167074
rect 267096 167010 267148 167016
rect 266452 159996 266504 160002
rect 266452 159938 266504 159944
rect 266360 144900 266412 144906
rect 266360 144842 266412 144848
rect 267004 136808 267056 136814
rect 267004 136750 267056 136756
rect 265900 136536 265952 136542
rect 265900 136478 265952 136484
rect 265808 120080 265860 120086
rect 265808 120022 265860 120028
rect 267016 65618 267044 136750
rect 267108 128246 267136 167010
rect 267200 130966 267228 169730
rect 267752 147626 267780 187138
rect 267844 164218 267872 203730
rect 267924 177540 267976 177546
rect 267924 177482 267976 177488
rect 267832 164212 267884 164218
rect 267832 164154 267884 164160
rect 267936 154426 267964 177482
rect 267924 154420 267976 154426
rect 267924 154362 267976 154368
rect 267740 147620 267792 147626
rect 267740 147562 267792 147568
rect 267188 130960 267240 130966
rect 267188 130902 267240 130908
rect 267096 128240 267148 128246
rect 267096 128182 267148 128188
rect 267096 107908 267148 107914
rect 267096 107850 267148 107856
rect 267004 65612 267056 65618
rect 267004 65554 267056 65560
rect 267108 61470 267136 107850
rect 267832 84856 267884 84862
rect 267832 84798 267884 84804
rect 267096 61464 267148 61470
rect 267096 61406 267148 61412
rect 265716 11824 265768 11830
rect 265716 11766 265768 11772
rect 267844 6914 267872 84798
rect 267752 6886 267872 6914
rect 266544 6384 266596 6390
rect 266544 6326 266596 6332
rect 265624 4956 265676 4962
rect 265624 4898 265676 4904
rect 266556 480 266584 6326
rect 267752 480 267780 6886
rect 268396 3670 268424 227054
rect 273260 222896 273312 222902
rect 273260 222838 273312 222844
rect 269120 218952 269172 218958
rect 269120 218894 269172 218900
rect 268476 162920 268528 162926
rect 268476 162862 268528 162868
rect 268488 124098 268516 162862
rect 269132 155242 269160 218894
rect 270592 214872 270644 214878
rect 270592 214814 270644 214820
rect 269212 192500 269264 192506
rect 269212 192442 269264 192448
rect 269224 160070 269252 192442
rect 269304 188420 269356 188426
rect 269304 188362 269356 188368
rect 269212 160064 269264 160070
rect 269212 160006 269264 160012
rect 269316 157282 269344 188362
rect 270500 180260 270552 180266
rect 270500 180202 270552 180208
rect 269764 172644 269816 172650
rect 269764 172586 269816 172592
rect 269304 157276 269356 157282
rect 269304 157218 269356 157224
rect 269120 155236 269172 155242
rect 269120 155178 269172 155184
rect 269776 135182 269804 172586
rect 269856 156052 269908 156058
rect 269856 155994 269908 156000
rect 269868 142866 269896 155994
rect 269948 153332 270000 153338
rect 269948 153274 270000 153280
rect 269856 142860 269908 142866
rect 269856 142802 269908 142808
rect 269960 141409 269988 153274
rect 269946 141400 270002 141409
rect 269946 141335 270002 141344
rect 269764 135176 269816 135182
rect 269764 135118 269816 135124
rect 269948 134564 270000 134570
rect 269948 134506 270000 134512
rect 269856 128376 269908 128382
rect 269856 128318 269908 128324
rect 268476 124092 268528 124098
rect 268476 124034 268528 124040
rect 269764 118720 269816 118726
rect 269764 118662 269816 118668
rect 268476 114572 268528 114578
rect 268476 114514 268528 114520
rect 268488 47666 268516 114514
rect 268476 47660 268528 47666
rect 268476 47602 268528 47608
rect 269776 29714 269804 118662
rect 269868 43450 269896 128318
rect 269960 100570 269988 134506
rect 269948 100564 270000 100570
rect 269948 100506 270000 100512
rect 269856 43444 269908 43450
rect 269856 43386 269908 43392
rect 269764 29708 269816 29714
rect 269764 29650 269816 29656
rect 268844 4140 268896 4146
rect 268844 4082 268896 4088
rect 268384 3664 268436 3670
rect 268384 3606 268436 3612
rect 268856 480 268884 4082
rect 270512 3534 270540 180202
rect 270604 162858 270632 214814
rect 272064 211948 272116 211954
rect 272064 211890 272116 211896
rect 270684 206576 270736 206582
rect 270684 206518 270736 206524
rect 270696 165578 270724 206518
rect 271880 203720 271932 203726
rect 271880 203662 271932 203668
rect 271144 174004 271196 174010
rect 271144 173946 271196 173952
rect 270684 165572 270736 165578
rect 270684 165514 270736 165520
rect 270592 162852 270644 162858
rect 270592 162794 270644 162800
rect 271156 138786 271184 173946
rect 271236 164348 271288 164354
rect 271236 164290 271288 164296
rect 271144 138780 271196 138786
rect 271144 138722 271196 138728
rect 271144 127016 271196 127022
rect 271144 126958 271196 126964
rect 271156 36582 271184 126958
rect 271248 126954 271276 164290
rect 271328 142248 271380 142254
rect 271328 142190 271380 142196
rect 271236 126948 271288 126954
rect 271236 126890 271288 126896
rect 271236 109064 271288 109070
rect 271236 109006 271288 109012
rect 271248 55962 271276 109006
rect 271340 102134 271368 142190
rect 271328 102128 271380 102134
rect 271328 102070 271380 102076
rect 271236 55956 271288 55962
rect 271236 55898 271288 55904
rect 271144 36576 271196 36582
rect 271144 36518 271196 36524
rect 271892 16574 271920 203662
rect 271972 196716 272024 196722
rect 271972 196658 272024 196664
rect 271984 137970 272012 196658
rect 272076 154494 272104 211890
rect 272524 165708 272576 165714
rect 272524 165650 272576 165656
rect 272064 154488 272116 154494
rect 272064 154430 272116 154436
rect 272536 152590 272564 165650
rect 272524 152584 272576 152590
rect 272524 152526 272576 152532
rect 272616 147756 272668 147762
rect 272616 147698 272668 147704
rect 272524 138032 272576 138038
rect 272524 137974 272576 137980
rect 271972 137964 272024 137970
rect 271972 137906 272024 137912
rect 272536 58750 272564 137974
rect 272628 107642 272656 147698
rect 273272 146198 273300 222838
rect 273352 213308 273404 213314
rect 273352 213250 273404 213256
rect 273364 151638 273392 213250
rect 274640 206440 274692 206446
rect 274640 206382 274692 206388
rect 274088 174548 274140 174554
rect 274088 174490 274140 174496
rect 273904 169856 273956 169862
rect 273904 169798 273956 169804
rect 273352 151632 273404 151638
rect 273352 151574 273404 151580
rect 273260 146192 273312 146198
rect 273260 146134 273312 146140
rect 273916 131034 273944 169798
rect 273904 131028 273956 131034
rect 273904 130970 273956 130976
rect 273996 129804 274048 129810
rect 273996 129746 274048 129752
rect 273904 120148 273956 120154
rect 273904 120090 273956 120096
rect 272616 107636 272668 107642
rect 272616 107578 272668 107584
rect 272524 58744 272576 58750
rect 272524 58686 272576 58692
rect 273260 26988 273312 26994
rect 273260 26930 273312 26936
rect 271892 16546 272472 16574
rect 271236 3732 271288 3738
rect 271236 3674 271288 3680
rect 270500 3528 270552 3534
rect 270500 3470 270552 3476
rect 270040 3256 270092 3262
rect 270040 3198 270092 3204
rect 270052 480 270080 3198
rect 271248 480 271276 3674
rect 272444 480 272472 16546
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 26930
rect 273916 25566 273944 120090
rect 274008 37942 274036 129746
rect 274100 86970 274128 174490
rect 274180 150544 274232 150550
rect 274180 150486 274232 150492
rect 274192 110362 274220 150486
rect 274180 110356 274232 110362
rect 274180 110298 274232 110304
rect 274180 99408 274232 99414
rect 274180 99350 274232 99356
rect 274088 86964 274140 86970
rect 274088 86906 274140 86912
rect 274192 39370 274220 99350
rect 274180 39364 274232 39370
rect 274180 39306 274232 39312
rect 273996 37936 274048 37942
rect 273996 37878 274048 37884
rect 273904 25560 273956 25566
rect 273904 25502 273956 25508
rect 274652 16574 274680 206382
rect 274824 190120 274876 190126
rect 274824 190062 274876 190068
rect 274732 184476 274784 184482
rect 274732 184418 274784 184424
rect 274744 150414 274772 184418
rect 274836 157350 274864 190062
rect 274824 157344 274876 157350
rect 274824 157286 274876 157292
rect 274732 150408 274784 150414
rect 274732 150350 274784 150356
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 275296 3602 275324 235311
rect 277412 224942 277440 240094
rect 278780 236700 278832 236706
rect 278780 236642 278832 236648
rect 277400 224936 277452 224942
rect 277400 224878 277452 224884
rect 278044 220108 278096 220114
rect 278044 220050 278096 220056
rect 277400 209092 277452 209098
rect 277400 209034 277452 209040
rect 276112 198144 276164 198150
rect 276112 198086 276164 198092
rect 276020 196648 276072 196654
rect 276020 196590 276072 196596
rect 275560 151836 275612 151842
rect 275560 151778 275612 151784
rect 275468 140820 275520 140826
rect 275468 140762 275520 140768
rect 275376 110492 275428 110498
rect 275376 110434 275428 110440
rect 275388 51814 275416 110434
rect 275480 100638 275508 140762
rect 275572 111790 275600 151778
rect 276032 146266 276060 196590
rect 276124 155922 276152 198086
rect 276112 155916 276164 155922
rect 276112 155858 276164 155864
rect 276756 154692 276808 154698
rect 276756 154634 276808 154640
rect 276664 149184 276716 149190
rect 276664 149126 276716 149132
rect 276020 146260 276072 146266
rect 276020 146202 276072 146208
rect 276020 126336 276072 126342
rect 276020 126278 276072 126284
rect 275560 111784 275612 111790
rect 275560 111726 275612 111732
rect 275468 100632 275520 100638
rect 275468 100574 275520 100580
rect 275376 51808 275428 51814
rect 275376 51750 275428 51756
rect 276032 16574 276060 126278
rect 276676 108934 276704 149126
rect 276768 114442 276796 154634
rect 277412 154562 277440 209034
rect 277400 154556 277452 154562
rect 277400 154498 277452 154504
rect 276756 114436 276808 114442
rect 276756 114378 276808 114384
rect 276664 108928 276716 108934
rect 276664 108870 276716 108876
rect 276664 106412 276716 106418
rect 276664 106354 276716 106360
rect 276676 31074 276704 106354
rect 276664 31068 276716 31074
rect 276664 31010 276716 31016
rect 276032 16546 276704 16574
rect 276020 6316 276072 6322
rect 276020 6258 276072 6264
rect 275284 3596 275336 3602
rect 275284 3538 275336 3544
rect 276032 480 276060 6258
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278056 3602 278084 220050
rect 278136 164416 278188 164422
rect 278136 164358 278188 164364
rect 278148 135998 278176 164358
rect 278412 156664 278464 156670
rect 278412 156606 278464 156612
rect 278136 135992 278188 135998
rect 278136 135934 278188 135940
rect 278320 135312 278372 135318
rect 278320 135254 278372 135260
rect 278228 129872 278280 129878
rect 278228 129814 278280 129820
rect 278136 116068 278188 116074
rect 278136 116010 278188 116016
rect 278148 4826 278176 116010
rect 278240 39438 278268 129814
rect 278332 66978 278360 135254
rect 278424 117298 278452 156606
rect 278412 117292 278464 117298
rect 278412 117234 278464 117240
rect 278320 66972 278372 66978
rect 278320 66914 278372 66920
rect 278228 39432 278280 39438
rect 278228 39374 278280 39380
rect 278792 16574 278820 236642
rect 278884 231742 278912 240094
rect 278872 231736 278924 231742
rect 278872 231678 278924 231684
rect 280160 215960 280212 215966
rect 280160 215902 280212 215908
rect 278964 205012 279016 205018
rect 278964 204954 279016 204960
rect 278872 202224 278924 202230
rect 278872 202166 278924 202172
rect 278884 139398 278912 202166
rect 278976 153202 279004 204954
rect 279424 168496 279476 168502
rect 279424 168438 279476 168444
rect 278964 153196 279016 153202
rect 278964 153138 279016 153144
rect 278872 139392 278924 139398
rect 278872 139334 278924 139340
rect 279436 131102 279464 168438
rect 280172 149054 280200 215902
rect 281552 203658 281580 240094
rect 284358 239850 284386 240108
rect 284312 239822 284386 239850
rect 285692 240094 286304 240122
rect 284312 237454 284340 239822
rect 283564 237448 283616 237454
rect 283564 237390 283616 237396
rect 284300 237448 284352 237454
rect 284300 237390 284352 237396
rect 282184 232552 282236 232558
rect 282184 232494 282236 232500
rect 281540 203652 281592 203658
rect 281540 203594 281592 203600
rect 281080 171216 281132 171222
rect 281080 171158 281132 171164
rect 280160 149048 280212 149054
rect 280160 148990 280212 148996
rect 279608 143676 279660 143682
rect 279608 143618 279660 143624
rect 279516 134088 279568 134094
rect 279516 134030 279568 134036
rect 279424 131096 279476 131102
rect 279424 131038 279476 131044
rect 279424 127084 279476 127090
rect 279424 127026 279476 127032
rect 278792 16546 279096 16574
rect 278136 4820 278188 4826
rect 278136 4762 278188 4768
rect 278318 4040 278374 4049
rect 278318 3975 278374 3984
rect 278044 3596 278096 3602
rect 278044 3538 278096 3544
rect 278332 480 278360 3975
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 279436 7614 279464 127026
rect 279528 72554 279556 134030
rect 279620 111110 279648 143618
rect 280896 139460 280948 139466
rect 280896 139402 280948 139408
rect 280804 133272 280856 133278
rect 280804 133214 280856 133220
rect 279608 111104 279660 111110
rect 279608 111046 279660 111052
rect 279516 72548 279568 72554
rect 279516 72490 279568 72496
rect 279424 7608 279476 7614
rect 279424 7550 279476 7556
rect 280816 3534 280844 133214
rect 280908 49026 280936 139402
rect 281092 133890 281120 171158
rect 281080 133884 281132 133890
rect 281080 133826 281132 133832
rect 280988 132524 281040 132530
rect 280988 132466 281040 132472
rect 281000 55894 281028 132466
rect 280988 55888 281040 55894
rect 280988 55830 281040 55836
rect 280896 49020 280948 49026
rect 280896 48962 280948 48968
rect 281908 9104 281960 9110
rect 281908 9046 281960 9052
rect 280804 3528 280856 3534
rect 280804 3470 280856 3476
rect 280712 3460 280764 3466
rect 280712 3402 280764 3408
rect 280724 480 280752 3402
rect 281920 480 281948 9046
rect 282196 3466 282224 232494
rect 282368 165776 282420 165782
rect 282368 165718 282420 165724
rect 282276 132592 282328 132598
rect 282276 132534 282328 132540
rect 282288 57322 282316 132534
rect 282380 128314 282408 165718
rect 282460 153876 282512 153882
rect 282460 153818 282512 153824
rect 282368 128308 282420 128314
rect 282368 128250 282420 128256
rect 282368 116136 282420 116142
rect 282368 116078 282420 116084
rect 282276 57316 282328 57322
rect 282276 57258 282328 57264
rect 282380 42090 282408 116078
rect 282472 115938 282500 153818
rect 282460 115932 282512 115938
rect 282460 115874 282512 115880
rect 283576 95946 283604 237390
rect 283656 220244 283708 220250
rect 283656 220186 283708 220192
rect 283668 178673 283696 220186
rect 283654 178664 283710 178673
rect 283654 178599 283710 178608
rect 283656 172712 283708 172718
rect 283656 172654 283708 172660
rect 283668 135250 283696 172654
rect 283748 160200 283800 160206
rect 283748 160142 283800 160148
rect 283656 135244 283708 135250
rect 283656 135186 283708 135192
rect 283656 121576 283708 121582
rect 283656 121518 283708 121524
rect 283564 95940 283616 95946
rect 283564 95882 283616 95888
rect 282368 42084 282420 42090
rect 282368 42026 282420 42032
rect 283668 19990 283696 121518
rect 283760 121378 283788 160142
rect 285220 154760 285272 154766
rect 285220 154702 285272 154708
rect 285128 151904 285180 151910
rect 285128 151846 285180 151852
rect 284944 146464 284996 146470
rect 284944 146406 284996 146412
rect 283840 131164 283892 131170
rect 283840 131106 283892 131112
rect 283748 121372 283800 121378
rect 283748 121314 283800 121320
rect 283748 110560 283800 110566
rect 283748 110502 283800 110508
rect 283656 19984 283708 19990
rect 283656 19926 283708 19932
rect 283760 18630 283788 110502
rect 283852 54534 283880 131106
rect 284956 123486 284984 146406
rect 285140 131782 285168 151846
rect 285128 131776 285180 131782
rect 285128 131718 285180 131724
rect 285036 131232 285088 131238
rect 285036 131174 285088 131180
rect 284944 123480 284996 123486
rect 284944 123422 284996 123428
rect 284944 113212 284996 113218
rect 284944 113154 284996 113160
rect 283840 54528 283892 54534
rect 283840 54470 283892 54476
rect 284956 29646 284984 113154
rect 285048 53106 285076 131174
rect 285128 122868 285180 122874
rect 285128 122810 285180 122816
rect 285140 75206 285168 122810
rect 285232 114510 285260 154702
rect 285220 114504 285272 114510
rect 285220 114446 285272 114452
rect 285128 75200 285180 75206
rect 285128 75142 285180 75148
rect 285036 53100 285088 53106
rect 285036 53042 285088 53048
rect 284944 29640 284996 29646
rect 284944 29582 284996 29588
rect 283748 18624 283800 18630
rect 283748 18566 283800 18572
rect 284300 6452 284352 6458
rect 284300 6394 284352 6400
rect 283104 3664 283156 3670
rect 283104 3606 283156 3612
rect 282184 3460 282236 3466
rect 282184 3402 282236 3408
rect 283116 480 283144 3606
rect 284312 480 284340 6394
rect 285692 3482 285720 240094
rect 287702 240071 287758 240080
rect 287716 227730 287744 240071
rect 288222 239850 288250 240108
rect 288176 239822 288250 239850
rect 290476 240094 290812 240122
rect 288176 238610 288204 239822
rect 288164 238604 288216 238610
rect 288164 238546 288216 238552
rect 288176 233238 288204 238546
rect 290476 237182 290504 240094
rect 291936 237448 291988 237454
rect 291936 237390 291988 237396
rect 290464 237176 290516 237182
rect 290464 237118 290516 237124
rect 288164 233232 288216 233238
rect 288164 233174 288216 233180
rect 287704 227724 287756 227730
rect 287704 227666 287756 227672
rect 290476 226302 290504 237118
rect 290464 226296 290516 226302
rect 290464 226238 290516 226244
rect 287796 222964 287848 222970
rect 287796 222906 287848 222912
rect 287704 206644 287756 206650
rect 287704 206586 287756 206592
rect 286324 128444 286376 128450
rect 286324 128386 286376 128392
rect 285772 83564 285824 83570
rect 285772 83506 285824 83512
rect 285784 16574 285812 83506
rect 286336 33794 286364 128386
rect 286324 33788 286376 33794
rect 286324 33730 286376 33736
rect 285784 16546 286640 16574
rect 285416 3454 285720 3482
rect 285416 480 285444 3454
rect 286612 480 286640 16546
rect 287336 10396 287388 10402
rect 287336 10338 287388 10344
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 10338
rect 287716 3534 287744 206586
rect 287808 177342 287836 222906
rect 289820 211200 289872 211206
rect 289820 211142 289872 211148
rect 289084 210452 289136 210458
rect 289084 210394 289136 210400
rect 289096 181626 289124 210394
rect 289084 181620 289136 181626
rect 289084 181562 289136 181568
rect 289084 178084 289136 178090
rect 289084 178026 289136 178032
rect 287796 177336 287848 177342
rect 287796 177278 287848 177284
rect 287980 174072 288032 174078
rect 287980 174014 288032 174020
rect 287888 168564 287940 168570
rect 287888 168506 287940 168512
rect 287900 129742 287928 168506
rect 287888 129736 287940 129742
rect 287888 129678 287940 129684
rect 287796 128512 287848 128518
rect 287796 128454 287848 128460
rect 287808 46306 287836 128454
rect 287888 122936 287940 122942
rect 287888 122878 287940 122884
rect 287796 46300 287848 46306
rect 287796 46242 287848 46248
rect 287900 43518 287928 122878
rect 287992 104174 288020 174014
rect 287980 104168 288032 104174
rect 287980 104110 288032 104116
rect 289096 101454 289124 178026
rect 289728 177404 289780 177410
rect 289728 177346 289780 177352
rect 289360 140888 289412 140894
rect 289360 140830 289412 140836
rect 289176 125724 289228 125730
rect 289176 125666 289228 125672
rect 289084 101448 289136 101454
rect 289084 101390 289136 101396
rect 289084 96824 289136 96830
rect 289084 96766 289136 96772
rect 287888 43512 287940 43518
rect 287888 43454 287940 43460
rect 289096 8974 289124 96766
rect 289188 40730 289216 125666
rect 289372 100706 289400 140830
rect 289360 100700 289412 100706
rect 289360 100642 289412 100648
rect 289268 99476 289320 99482
rect 289268 99418 289320 99424
rect 289280 46238 289308 99418
rect 289268 46232 289320 46238
rect 289268 46174 289320 46180
rect 289176 40724 289228 40730
rect 289176 40666 289228 40672
rect 289084 8968 289136 8974
rect 289084 8910 289136 8916
rect 289740 3602 289768 177346
rect 288992 3596 289044 3602
rect 288992 3538 289044 3544
rect 289728 3596 289780 3602
rect 289728 3538 289780 3544
rect 287704 3528 287756 3534
rect 287704 3470 287756 3476
rect 289004 480 289032 3538
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 211142
rect 291844 163532 291896 163538
rect 291844 163474 291896 163480
rect 290648 162988 290700 162994
rect 290648 162930 290700 162936
rect 290556 138100 290608 138106
rect 290556 138042 290608 138048
rect 290464 123004 290516 123010
rect 290464 122946 290516 122952
rect 290476 31142 290504 122946
rect 290568 62830 290596 138042
rect 290660 124166 290688 162930
rect 290648 124160 290700 124166
rect 290648 124102 290700 124108
rect 290556 62824 290608 62830
rect 290556 62766 290608 62772
rect 290464 31136 290516 31142
rect 290464 31078 290516 31084
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 291396 480 291424 3470
rect 291856 3466 291884 163474
rect 291948 86290 291976 237390
rect 292040 126342 292068 240586
rect 292592 240094 292744 240122
rect 292592 237454 292620 240094
rect 292670 239184 292726 239193
rect 292670 239119 292672 239128
rect 292724 239119 292726 239128
rect 292672 239090 292724 239096
rect 292580 237448 292632 237454
rect 292580 237390 292632 237396
rect 292028 126336 292080 126342
rect 292028 126278 292080 126284
rect 292028 117360 292080 117366
rect 292028 117302 292080 117308
rect 291936 86284 291988 86290
rect 291936 86226 291988 86232
rect 292040 21486 292068 117302
rect 292120 100836 292172 100842
rect 292120 100778 292172 100784
rect 292028 21480 292080 21486
rect 292028 21422 292080 21428
rect 292132 11762 292160 100778
rect 293052 83570 293080 346967
rect 293144 314265 293172 354719
rect 293236 334665 293264 368863
rect 293972 357377 294000 387806
rect 294052 381608 294104 381614
rect 294052 381550 294104 381556
rect 293958 357368 294014 357377
rect 293958 357303 294014 357312
rect 293316 354544 293368 354550
rect 293314 354512 293316 354521
rect 293368 354512 293370 354521
rect 293314 354447 293370 354456
rect 293958 352336 294014 352345
rect 293958 352271 294014 352280
rect 293222 334656 293278 334665
rect 293222 334591 293278 334600
rect 293130 314256 293186 314265
rect 293130 314191 293186 314200
rect 293866 314256 293922 314265
rect 293866 314191 293922 314200
rect 293880 313342 293908 314191
rect 293868 313336 293920 313342
rect 293868 313278 293920 313284
rect 293130 287736 293186 287745
rect 293130 287671 293186 287680
rect 293144 117978 293172 287671
rect 293222 259176 293278 259185
rect 293222 259111 293278 259120
rect 293236 206446 293264 259111
rect 293314 241224 293370 241233
rect 293314 241159 293370 241168
rect 293328 240650 293356 241159
rect 293316 240644 293368 240650
rect 293316 240586 293368 240592
rect 293224 206440 293276 206446
rect 293224 206382 293276 206388
rect 293224 118788 293276 118794
rect 293224 118730 293276 118736
rect 293132 117972 293184 117978
rect 293132 117914 293184 117920
rect 293040 83564 293092 83570
rect 293040 83506 293092 83512
rect 293236 14482 293264 118730
rect 293316 103556 293368 103562
rect 293316 103498 293368 103504
rect 293328 33862 293356 103498
rect 293972 102814 294000 352271
rect 294064 331945 294092 381550
rect 295616 374060 295668 374066
rect 295616 374002 295668 374008
rect 295524 373312 295576 373318
rect 295524 373254 295576 373260
rect 295340 371884 295392 371890
rect 295340 371826 295392 371832
rect 294144 369164 294196 369170
rect 294144 369106 294196 369112
rect 294156 336705 294184 369106
rect 294236 356244 294288 356250
rect 294236 356186 294288 356192
rect 294142 336696 294198 336705
rect 294142 336631 294198 336640
rect 294050 331936 294106 331945
rect 294050 331871 294106 331880
rect 294050 325816 294106 325825
rect 294050 325751 294106 325760
rect 294064 203726 294092 325751
rect 294142 312216 294198 312225
rect 294142 312151 294198 312160
rect 294156 229090 294184 312151
rect 294248 309097 294276 356186
rect 295352 310706 295380 371826
rect 295432 362364 295484 362370
rect 295432 362306 295484 362312
rect 295444 325694 295472 362306
rect 295536 361690 295564 373254
rect 295524 361684 295576 361690
rect 295524 361626 295576 361632
rect 295536 327865 295564 361626
rect 295628 345710 295656 374002
rect 295616 345704 295668 345710
rect 295616 345646 295668 345652
rect 295628 345545 295656 345646
rect 295614 345536 295670 345545
rect 295614 345471 295670 345480
rect 296732 343670 296760 512586
rect 297376 400110 297404 702714
rect 299492 594114 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 299480 594108 299532 594114
rect 299480 594050 299532 594056
rect 331232 588606 331260 702986
rect 348804 697610 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 697604 348844 697610
rect 348792 697546 348844 697552
rect 363604 696992 363656 696998
rect 363604 696934 363656 696940
rect 331220 588600 331272 588606
rect 331220 588542 331272 588548
rect 336740 582412 336792 582418
rect 336740 582354 336792 582360
rect 335360 575544 335412 575550
rect 335360 575486 335412 575492
rect 332600 565888 332652 565894
rect 332600 565830 332652 565836
rect 314660 556232 314712 556238
rect 314660 556174 314712 556180
rect 313280 536104 313332 536110
rect 313280 536046 313332 536052
rect 300860 505776 300912 505782
rect 300860 505718 300912 505724
rect 299480 472660 299532 472666
rect 299480 472602 299532 472608
rect 299492 472054 299520 472602
rect 299480 472048 299532 472054
rect 299480 471990 299532 471996
rect 298192 411324 298244 411330
rect 298192 411266 298244 411272
rect 296812 400104 296864 400110
rect 296812 400046 296864 400052
rect 297364 400104 297416 400110
rect 297364 400046 297416 400052
rect 296076 343664 296128 343670
rect 296076 343606 296128 343612
rect 296720 343664 296772 343670
rect 296720 343606 296772 343612
rect 295614 340776 295670 340785
rect 295614 340711 295670 340720
rect 295628 339522 295656 340711
rect 295616 339516 295668 339522
rect 295616 339458 295668 339464
rect 295616 339176 295668 339182
rect 295616 339118 295668 339124
rect 295628 338745 295656 339118
rect 295614 338736 295670 338745
rect 295614 338671 295670 338680
rect 295522 327856 295578 327865
rect 295522 327791 295578 327800
rect 295536 327758 295564 327791
rect 295524 327752 295576 327758
rect 295524 327694 295576 327700
rect 295444 325666 295656 325694
rect 295430 321056 295486 321065
rect 295430 320991 295486 321000
rect 295444 320210 295472 320991
rect 295432 320204 295484 320210
rect 295432 320146 295484 320152
rect 295430 319016 295486 319025
rect 295430 318951 295486 318960
rect 295444 318850 295472 318951
rect 295432 318844 295484 318850
rect 295432 318786 295484 318792
rect 295432 317416 295484 317422
rect 295432 317358 295484 317364
rect 295444 316985 295472 317358
rect 295430 316976 295486 316985
rect 295430 316911 295486 316920
rect 295352 310678 295564 310706
rect 295340 310480 295392 310486
rect 295340 310422 295392 310428
rect 295352 310185 295380 310422
rect 295338 310176 295394 310185
rect 295338 310111 295394 310120
rect 294234 309088 294290 309097
rect 294234 309023 294290 309032
rect 295536 308446 295564 310678
rect 295524 308440 295576 308446
rect 295524 308382 295576 308388
rect 295536 308145 295564 308382
rect 295522 308136 295578 308145
rect 295522 308071 295578 308080
rect 295338 301336 295394 301345
rect 295338 301271 295394 301280
rect 295352 300898 295380 301271
rect 295340 300892 295392 300898
rect 295340 300834 295392 300840
rect 295338 299296 295394 299305
rect 295338 299231 295394 299240
rect 295352 294658 295380 299231
rect 295628 296714 295656 325666
rect 295260 294630 295380 294658
rect 295444 296686 295656 296714
rect 295260 293842 295288 294630
rect 295338 294536 295394 294545
rect 295338 294471 295394 294480
rect 295352 294030 295380 294471
rect 295340 294024 295392 294030
rect 295340 293966 295392 293972
rect 295260 293814 295380 293842
rect 294234 268016 294290 268025
rect 294234 267951 294290 267960
rect 294248 236706 294276 267951
rect 294236 236700 294288 236706
rect 294236 236642 294288 236648
rect 294144 229084 294196 229090
rect 294144 229026 294196 229032
rect 294052 203720 294104 203726
rect 294052 203662 294104 203668
rect 294604 167748 294656 167754
rect 294604 167690 294656 167696
rect 294616 136610 294644 167690
rect 294604 136604 294656 136610
rect 294604 136546 294656 136552
rect 294696 135380 294748 135386
rect 294696 135322 294748 135328
rect 294604 113280 294656 113286
rect 294604 113222 294656 113228
rect 293960 102808 294012 102814
rect 293960 102750 294012 102756
rect 293408 98184 293460 98190
rect 293408 98126 293460 98132
rect 293420 73846 293448 98126
rect 293408 73840 293460 73846
rect 293408 73782 293460 73788
rect 294616 35222 294644 113222
rect 294708 68406 294736 135322
rect 294788 127628 294840 127634
rect 294788 127570 294840 127576
rect 294800 104854 294828 127570
rect 295352 105602 295380 293814
rect 295444 287054 295472 296686
rect 295522 296576 295578 296585
rect 295522 296511 295578 296520
rect 295536 295390 295564 296511
rect 295524 295384 295576 295390
rect 295524 295326 295576 295332
rect 295614 292496 295670 292505
rect 295614 292431 295670 292440
rect 295628 291242 295656 292431
rect 295616 291236 295668 291242
rect 295616 291178 295668 291184
rect 295524 291168 295576 291174
rect 295524 291110 295576 291116
rect 295536 290465 295564 291110
rect 295522 290456 295578 290465
rect 295522 290391 295578 290400
rect 295444 287026 295564 287054
rect 295432 285728 295484 285734
rect 295430 285696 295432 285705
rect 295484 285696 295486 285705
rect 295430 285631 295486 285640
rect 295430 283656 295486 283665
rect 295536 283642 295564 287026
rect 295486 283614 295564 283642
rect 295430 283591 295432 283600
rect 295484 283591 295486 283600
rect 295432 283562 295484 283568
rect 295430 281616 295486 281625
rect 295430 281551 295432 281560
rect 295484 281551 295486 281560
rect 295432 281522 295484 281528
rect 295430 278896 295486 278905
rect 295430 278831 295432 278840
rect 295484 278831 295486 278840
rect 295432 278802 295484 278808
rect 295430 276856 295486 276865
rect 295430 276791 295486 276800
rect 295444 276078 295472 276791
rect 295432 276072 295484 276078
rect 295432 276014 295484 276020
rect 295430 274816 295486 274825
rect 295430 274751 295486 274760
rect 295444 274718 295472 274751
rect 295432 274712 295484 274718
rect 295432 274654 295484 274660
rect 295430 272776 295486 272785
rect 295430 272711 295432 272720
rect 295484 272711 295486 272720
rect 295432 272682 295484 272688
rect 295430 270056 295486 270065
rect 295430 269991 295486 270000
rect 295444 269142 295472 269991
rect 295432 269136 295484 269142
rect 295432 269078 295484 269084
rect 295430 265976 295486 265985
rect 295430 265911 295486 265920
rect 295444 264994 295472 265911
rect 295432 264988 295484 264994
rect 295432 264930 295484 264936
rect 295522 263936 295578 263945
rect 295522 263871 295578 263880
rect 295430 261216 295486 261225
rect 295430 261151 295486 261160
rect 295444 260914 295472 261151
rect 295432 260908 295484 260914
rect 295432 260850 295484 260856
rect 295536 258074 295564 263871
rect 295444 258046 295564 258074
rect 295340 105596 295392 105602
rect 295340 105538 295392 105544
rect 294788 104848 294840 104854
rect 294788 104790 294840 104796
rect 294880 103624 294932 103630
rect 294880 103566 294932 103572
rect 294788 102264 294840 102270
rect 294788 102206 294840 102212
rect 294696 68400 294748 68406
rect 294696 68342 294748 68348
rect 294800 44878 294828 102206
rect 294892 69698 294920 103566
rect 295444 84930 295472 258046
rect 295522 255096 295578 255105
rect 295522 255031 295578 255040
rect 295536 253978 295564 255031
rect 295524 253972 295576 253978
rect 295524 253914 295576 253920
rect 295522 252376 295578 252385
rect 295522 252311 295578 252320
rect 295536 251870 295564 252311
rect 295524 251864 295576 251870
rect 295524 251806 295576 251812
rect 295522 250336 295578 250345
rect 295522 250271 295578 250280
rect 295536 249830 295564 250271
rect 295524 249824 295576 249830
rect 295524 249766 295576 249772
rect 295522 246256 295578 246265
rect 295522 246191 295578 246200
rect 295536 245682 295564 246191
rect 295524 245676 295576 245682
rect 295524 245618 295576 245624
rect 295536 233102 295564 245618
rect 296088 238542 296116 343606
rect 296626 343496 296682 343505
rect 296824 343482 296852 400046
rect 296904 364472 296956 364478
rect 296904 364414 296956 364420
rect 296682 343454 296852 343482
rect 296626 343431 296682 343440
rect 296626 323096 296682 323105
rect 296682 323054 296760 323082
rect 296626 323031 296682 323040
rect 296076 238536 296128 238542
rect 296076 238478 296128 238484
rect 295524 233096 295576 233102
rect 295524 233038 295576 233044
rect 296732 211206 296760 323054
rect 296824 233170 296852 343454
rect 296916 329905 296944 364414
rect 298100 357604 298152 357610
rect 298100 357546 298152 357552
rect 297364 355020 297416 355026
rect 297364 354962 297416 354968
rect 296902 329896 296958 329905
rect 296902 329831 296958 329840
rect 297376 299470 297404 354962
rect 297364 299464 297416 299470
rect 297364 299406 297416 299412
rect 297364 278860 297416 278866
rect 297364 278802 297416 278808
rect 296902 243536 296958 243545
rect 296902 243471 296958 243480
rect 296916 242962 296944 243471
rect 296904 242956 296956 242962
rect 296904 242898 296956 242904
rect 296916 237318 296944 242898
rect 296904 237312 296956 237318
rect 296904 237254 296956 237260
rect 296812 233164 296864 233170
rect 296812 233106 296864 233112
rect 296720 211200 296772 211206
rect 296720 211142 296772 211148
rect 296076 157548 296128 157554
rect 296076 157490 296128 157496
rect 295984 134020 296036 134026
rect 295984 133962 296036 133968
rect 295432 84924 295484 84930
rect 295432 84866 295484 84872
rect 294880 69692 294932 69698
rect 294880 69634 294932 69640
rect 294788 44872 294840 44878
rect 294788 44814 294840 44820
rect 294604 35216 294656 35222
rect 294604 35158 294656 35164
rect 293316 33856 293368 33862
rect 293316 33798 293368 33804
rect 293224 14476 293276 14482
rect 293224 14418 293276 14424
rect 294880 11892 294932 11898
rect 294880 11834 294932 11840
rect 292120 11756 292172 11762
rect 292120 11698 292172 11704
rect 292580 6248 292632 6254
rect 292580 6190 292632 6196
rect 291844 3460 291896 3466
rect 291844 3402 291896 3408
rect 292592 480 292620 6190
rect 293684 3596 293736 3602
rect 293684 3538 293736 3544
rect 293696 480 293724 3538
rect 294892 480 294920 11834
rect 295996 10334 296024 133962
rect 296088 118658 296116 157490
rect 296076 118652 296128 118658
rect 296076 118594 296128 118600
rect 296076 105052 296128 105058
rect 296076 104994 296128 105000
rect 296088 66910 296116 104994
rect 296168 102332 296220 102338
rect 296168 102274 296220 102280
rect 296180 72486 296208 102274
rect 296168 72480 296220 72486
rect 296168 72422 296220 72428
rect 296076 66904 296128 66910
rect 296076 66846 296128 66852
rect 297376 27606 297404 278802
rect 297548 138168 297600 138174
rect 297548 138110 297600 138116
rect 297456 117428 297508 117434
rect 297456 117370 297508 117376
rect 297364 27600 297416 27606
rect 297364 27542 297416 27548
rect 296720 25628 296772 25634
rect 296720 25570 296772 25576
rect 296732 16574 296760 25570
rect 296732 16546 297312 16574
rect 295984 10328 296036 10334
rect 295984 10270 296036 10276
rect 296074 4040 296130 4049
rect 296074 3975 296130 3984
rect 296088 480 296116 3975
rect 297284 480 297312 16546
rect 297468 2106 297496 117370
rect 297560 71194 297588 138110
rect 298112 133278 298140 357546
rect 298204 238882 298232 411266
rect 298284 361616 298336 361622
rect 298284 361558 298336 361564
rect 298296 339182 298324 361558
rect 298284 339176 298336 339182
rect 298284 339118 298336 339124
rect 298284 272740 298336 272746
rect 298284 272682 298336 272688
rect 298296 241466 298324 272682
rect 298376 251864 298428 251870
rect 298376 251806 298428 251812
rect 298284 241460 298336 241466
rect 298284 241402 298336 241408
rect 298192 238876 298244 238882
rect 298192 238818 298244 238824
rect 298388 231810 298416 251806
rect 299492 237114 299520 471990
rect 299572 402348 299624 402354
rect 299572 402290 299624 402296
rect 299584 238746 299612 402290
rect 300124 354952 300176 354958
rect 300124 354894 300176 354900
rect 300136 313274 300164 354894
rect 300124 313268 300176 313274
rect 300124 313210 300176 313216
rect 300124 295384 300176 295390
rect 300124 295326 300176 295332
rect 299572 238740 299624 238746
rect 299572 238682 299624 238688
rect 299480 237108 299532 237114
rect 299480 237050 299532 237056
rect 298376 231804 298428 231810
rect 298376 231746 298428 231752
rect 298744 161560 298796 161566
rect 298744 161502 298796 161508
rect 298100 133272 298152 133278
rect 298100 133214 298152 133220
rect 298756 122806 298784 161502
rect 299020 145036 299072 145042
rect 299020 144978 299072 144984
rect 298744 122800 298796 122806
rect 298744 122742 298796 122748
rect 298928 120216 298980 120222
rect 298928 120158 298980 120164
rect 297640 114640 297692 114646
rect 297640 114582 297692 114588
rect 297548 71188 297600 71194
rect 297548 71130 297600 71136
rect 297652 64190 297680 114582
rect 298836 111920 298888 111926
rect 298836 111862 298888 111868
rect 298744 104984 298796 104990
rect 298744 104926 298796 104932
rect 297640 64184 297692 64190
rect 297640 64126 297692 64132
rect 298756 7682 298784 104926
rect 298848 22778 298876 111862
rect 298940 50454 298968 120158
rect 299032 112470 299060 144978
rect 299112 144220 299164 144226
rect 299112 144162 299164 144168
rect 299020 112464 299072 112470
rect 299020 112406 299072 112412
rect 299020 109132 299072 109138
rect 299020 109074 299072 109080
rect 299032 54602 299060 109074
rect 299124 106282 299152 144162
rect 299112 106276 299164 106282
rect 299112 106218 299164 106224
rect 300136 87718 300164 295326
rect 300872 237182 300900 505718
rect 305000 496868 305052 496874
rect 305000 496810 305052 496816
rect 301044 365016 301096 365022
rect 301044 364958 301096 364964
rect 300952 354884 301004 354890
rect 300952 354826 301004 354832
rect 300860 237176 300912 237182
rect 300860 237118 300912 237124
rect 300964 138718 300992 354826
rect 301056 291174 301084 364958
rect 302332 360324 302384 360330
rect 302332 360266 302384 360272
rect 302240 358896 302292 358902
rect 302240 358838 302292 358844
rect 301228 291236 301280 291242
rect 301228 291178 301280 291184
rect 301044 291168 301096 291174
rect 301044 291110 301096 291116
rect 301136 274712 301188 274718
rect 301136 274654 301188 274660
rect 301148 241097 301176 274654
rect 301134 241088 301190 241097
rect 301134 241023 301190 241032
rect 301240 239902 301268 291178
rect 301228 239896 301280 239902
rect 301228 239838 301280 239844
rect 301504 158840 301556 158846
rect 301504 158782 301556 158788
rect 300952 138712 301004 138718
rect 300952 138654 301004 138660
rect 301516 124914 301544 158782
rect 301688 142316 301740 142322
rect 301688 142258 301740 142264
rect 301596 132660 301648 132666
rect 301596 132602 301648 132608
rect 301504 124908 301556 124914
rect 301504 124850 301556 124856
rect 300216 121644 300268 121650
rect 300216 121586 300268 121592
rect 300124 87712 300176 87718
rect 300124 87654 300176 87660
rect 299020 54596 299072 54602
rect 299020 54538 299072 54544
rect 298928 50448 298980 50454
rect 298928 50390 298980 50396
rect 300228 32434 300256 121586
rect 301504 118856 301556 118862
rect 301504 118798 301556 118804
rect 300308 111988 300360 111994
rect 300308 111930 300360 111936
rect 300320 42158 300348 111930
rect 300400 107772 300452 107778
rect 300400 107714 300452 107720
rect 300412 58682 300440 107714
rect 300400 58676 300452 58682
rect 300400 58618 300452 58624
rect 300308 42152 300360 42158
rect 300308 42094 300360 42100
rect 300216 32428 300268 32434
rect 300216 32370 300268 32376
rect 299480 27600 299532 27606
rect 299480 27542 299532 27548
rect 298836 22772 298888 22778
rect 298836 22714 298888 22720
rect 298744 7676 298796 7682
rect 298744 7618 298796 7624
rect 299492 3534 299520 27542
rect 299664 7744 299716 7750
rect 299664 7686 299716 7692
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 298468 3460 298520 3466
rect 298468 3402 298520 3408
rect 297456 2100 297508 2106
rect 297456 2042 297508 2048
rect 298480 480 298508 3402
rect 299676 480 299704 7686
rect 301516 6186 301544 118798
rect 301608 61402 301636 132602
rect 301700 110430 301728 142258
rect 302252 135930 302280 358838
rect 302344 317422 302372 360266
rect 304262 354648 304318 354657
rect 304262 354583 304318 354592
rect 302332 317416 302384 317422
rect 302332 317358 302384 317364
rect 302344 316742 302372 317358
rect 302332 316736 302384 316742
rect 302332 316678 302384 316684
rect 302332 308440 302384 308446
rect 302332 308382 302384 308388
rect 302344 235958 302372 308382
rect 302424 276072 302476 276078
rect 302424 276014 302476 276020
rect 302436 237250 302464 276014
rect 302424 237244 302476 237250
rect 302424 237186 302476 237192
rect 302332 235952 302384 235958
rect 302332 235894 302384 235900
rect 304276 216714 304304 354583
rect 305012 251870 305040 496810
rect 306380 433356 306432 433362
rect 306380 433298 306432 433304
rect 305184 357672 305236 357678
rect 305184 357614 305236 357620
rect 305092 354748 305144 354754
rect 305092 354690 305144 354696
rect 305000 251864 305052 251870
rect 305000 251806 305052 251812
rect 304264 216708 304316 216714
rect 304264 216650 304316 216656
rect 304264 169924 304316 169930
rect 304264 169866 304316 169872
rect 302976 160268 303028 160274
rect 302976 160210 303028 160216
rect 302240 135924 302292 135930
rect 302240 135866 302292 135872
rect 302884 135448 302936 135454
rect 302884 135390 302936 135396
rect 301780 124228 301832 124234
rect 301780 124170 301832 124176
rect 301688 110424 301740 110430
rect 301688 110366 301740 110372
rect 301688 106480 301740 106486
rect 301688 106422 301740 106428
rect 301596 61396 301648 61402
rect 301596 61338 301648 61344
rect 301700 36650 301728 106422
rect 301792 76634 301820 124170
rect 301780 76628 301832 76634
rect 301780 76570 301832 76576
rect 301688 36644 301740 36650
rect 301688 36586 301740 36592
rect 302896 17338 302924 135390
rect 302988 121446 303016 160210
rect 303160 149252 303212 149258
rect 303160 149194 303212 149200
rect 302976 121440 303028 121446
rect 302976 121382 303028 121388
rect 302976 117496 303028 117502
rect 302976 117438 303028 117444
rect 302988 24206 303016 117438
rect 303172 109002 303200 149194
rect 304276 132462 304304 169866
rect 304356 140956 304408 140962
rect 304356 140898 304408 140904
rect 304264 132456 304316 132462
rect 304264 132398 304316 132404
rect 304368 115161 304396 140898
rect 305104 130422 305132 354690
rect 305196 166326 305224 357614
rect 305276 356108 305328 356114
rect 305276 356050 305328 356056
rect 305288 310486 305316 356050
rect 305276 310480 305328 310486
rect 305276 310422 305328 310428
rect 305460 310480 305512 310486
rect 305460 310422 305512 310428
rect 305472 309806 305500 310422
rect 305460 309800 305512 309806
rect 305460 309742 305512 309748
rect 305276 300892 305328 300898
rect 305276 300834 305328 300840
rect 305288 231674 305316 300834
rect 306392 276078 306420 433298
rect 310612 408536 310664 408542
rect 310612 408478 310664 408484
rect 309140 402280 309192 402286
rect 309140 402222 309192 402228
rect 308404 357808 308456 357814
rect 308404 357750 308456 357756
rect 306472 356720 306524 356726
rect 306472 356662 306524 356668
rect 306380 276072 306432 276078
rect 306380 276014 306432 276020
rect 306484 235890 306512 356662
rect 307024 294024 307076 294030
rect 307024 293966 307076 293972
rect 306564 283620 306616 283626
rect 306564 283562 306616 283568
rect 306576 239970 306604 283562
rect 306564 239964 306616 239970
rect 306564 239906 306616 239912
rect 306472 235884 306524 235890
rect 306472 235826 306524 235832
rect 305276 231668 305328 231674
rect 305276 231610 305328 231616
rect 307036 175681 307064 293966
rect 307116 218816 307168 218822
rect 307116 218758 307168 218764
rect 307128 177313 307156 218758
rect 307114 177304 307170 177313
rect 307114 177239 307170 177248
rect 307022 175672 307078 175681
rect 307022 175607 307078 175616
rect 307574 175264 307630 175273
rect 307574 175199 307630 175208
rect 307022 174856 307078 174865
rect 307022 174791 307078 174800
rect 306930 172272 306986 172281
rect 306930 172207 306986 172216
rect 306944 171222 306972 172207
rect 306932 171216 306984 171222
rect 306932 171158 306984 171164
rect 307036 167754 307064 174791
rect 307298 174448 307354 174457
rect 307298 174383 307354 174392
rect 307312 174010 307340 174383
rect 307588 174078 307616 175199
rect 307576 174072 307628 174078
rect 307576 174014 307628 174020
rect 307666 174040 307722 174049
rect 307300 174004 307352 174010
rect 307666 173975 307722 173984
rect 307300 173946 307352 173952
rect 307680 173942 307708 173975
rect 307668 173936 307720 173942
rect 307668 173878 307720 173884
rect 307574 173632 307630 173641
rect 307574 173567 307630 173576
rect 307298 173224 307354 173233
rect 307298 173159 307354 173168
rect 307312 172650 307340 173159
rect 307588 172718 307616 173567
rect 307576 172712 307628 172718
rect 307576 172654 307628 172660
rect 307666 172680 307722 172689
rect 307300 172644 307352 172650
rect 307666 172615 307722 172624
rect 307300 172586 307352 172592
rect 307680 172582 307708 172615
rect 307668 172576 307720 172582
rect 307668 172518 307720 172524
rect 307482 171864 307538 171873
rect 307482 171799 307538 171808
rect 307496 171154 307524 171799
rect 307484 171148 307536 171154
rect 307484 171090 307536 171096
rect 307390 171048 307446 171057
rect 307390 170983 307446 170992
rect 307300 169856 307352 169862
rect 307298 169824 307300 169833
rect 307352 169824 307354 169833
rect 307298 169759 307354 169768
rect 307298 168464 307354 168473
rect 307298 168399 307300 168408
rect 307352 168399 307354 168408
rect 307300 168370 307352 168376
rect 307114 168056 307170 168065
rect 307114 167991 307170 168000
rect 307024 167748 307076 167754
rect 307024 167690 307076 167696
rect 306930 167648 306986 167657
rect 306930 167583 306986 167592
rect 306944 167074 306972 167583
rect 306932 167068 306984 167074
rect 306932 167010 306984 167016
rect 306930 166832 306986 166841
rect 306930 166767 306986 166776
rect 305184 166320 305236 166326
rect 305184 166262 305236 166268
rect 306944 165782 306972 166767
rect 306932 165776 306984 165782
rect 306932 165718 306984 165724
rect 305642 162888 305698 162897
rect 305642 162823 305698 162832
rect 305092 130416 305144 130422
rect 305092 130358 305144 130364
rect 305656 126274 305684 162823
rect 307022 161664 307078 161673
rect 307022 161599 307078 161608
rect 306746 161256 306802 161265
rect 306746 161191 306802 161200
rect 306760 160206 306788 161191
rect 306748 160200 306800 160206
rect 306748 160142 306800 160148
rect 306930 158672 306986 158681
rect 306930 158607 306986 158616
rect 306944 157486 306972 158607
rect 306932 157480 306984 157486
rect 306932 157422 306984 157428
rect 306746 157040 306802 157049
rect 306746 156975 306802 156984
rect 306760 155990 306788 156975
rect 306748 155984 306800 155990
rect 306748 155926 306800 155932
rect 306654 153232 306710 153241
rect 306654 153167 306710 153176
rect 306562 152280 306618 152289
rect 306562 152215 306618 152224
rect 306576 149734 306604 152215
rect 306668 151094 306696 153167
rect 306656 151088 306708 151094
rect 306656 151030 306708 151036
rect 306930 150240 306986 150249
rect 306930 150175 306986 150184
rect 306564 149728 306616 149734
rect 306564 149670 306616 149676
rect 306944 149190 306972 150175
rect 306932 149184 306984 149190
rect 306932 149126 306984 149132
rect 306746 147248 306802 147257
rect 306746 147183 306802 147192
rect 306760 146402 306788 147183
rect 306748 146396 306800 146402
rect 306748 146338 306800 146344
rect 307036 145586 307064 161599
rect 307128 160750 307156 167991
rect 307404 167686 307432 170983
rect 307482 170640 307538 170649
rect 307482 170575 307538 170584
rect 307496 169930 307524 170575
rect 307666 170232 307722 170241
rect 307666 170167 307722 170176
rect 307484 169924 307536 169930
rect 307484 169866 307536 169872
rect 307680 169794 307708 170167
rect 307668 169788 307720 169794
rect 307668 169730 307720 169736
rect 307574 169280 307630 169289
rect 307574 169215 307630 169224
rect 307588 168502 307616 169215
rect 307666 168872 307722 168881
rect 307666 168807 307722 168816
rect 307680 168570 307708 168807
rect 307668 168564 307720 168570
rect 307668 168506 307720 168512
rect 307576 168496 307628 168502
rect 307576 168438 307628 168444
rect 307392 167680 307444 167686
rect 307392 167622 307444 167628
rect 307206 167240 307262 167249
rect 307206 167175 307262 167184
rect 307220 162178 307248 167175
rect 307666 166424 307722 166433
rect 307666 166359 307722 166368
rect 307482 165880 307538 165889
rect 307482 165815 307538 165824
rect 307496 165714 307524 165815
rect 307484 165708 307536 165714
rect 307484 165650 307536 165656
rect 307680 165646 307708 166359
rect 307668 165640 307720 165646
rect 307668 165582 307720 165588
rect 307574 165472 307630 165481
rect 307574 165407 307630 165416
rect 307390 165064 307446 165073
rect 307390 164999 307446 165008
rect 307300 164280 307352 164286
rect 307298 164248 307300 164257
rect 307352 164248 307354 164257
rect 307298 164183 307354 164192
rect 307298 163432 307354 163441
rect 307298 163367 307354 163376
rect 307312 162994 307340 163367
rect 307300 162988 307352 162994
rect 307300 162930 307352 162936
rect 307208 162172 307260 162178
rect 307208 162114 307260 162120
rect 307116 160744 307168 160750
rect 307116 160686 307168 160692
rect 307404 159390 307432 164999
rect 307588 164354 307616 165407
rect 307666 164656 307722 164665
rect 307666 164591 307722 164600
rect 307680 164422 307708 164591
rect 307668 164416 307720 164422
rect 307668 164358 307720 164364
rect 307576 164348 307628 164354
rect 307576 164290 307628 164296
rect 307574 163840 307630 163849
rect 307574 163775 307630 163784
rect 307588 162897 307616 163775
rect 307666 163024 307722 163033
rect 307666 162959 307722 162968
rect 307680 162926 307708 162959
rect 307668 162920 307720 162926
rect 307574 162888 307630 162897
rect 307668 162862 307720 162868
rect 307574 162823 307630 162832
rect 307482 162480 307538 162489
rect 307482 162415 307538 162424
rect 307496 161566 307524 162415
rect 307666 162072 307722 162081
rect 307666 162007 307722 162016
rect 307484 161560 307536 161566
rect 307484 161502 307536 161508
rect 307680 161498 307708 162007
rect 307668 161492 307720 161498
rect 307668 161434 307720 161440
rect 307482 160848 307538 160857
rect 307482 160783 307538 160792
rect 307496 160138 307524 160783
rect 307666 160440 307722 160449
rect 307666 160375 307722 160384
rect 307680 160274 307708 160375
rect 307668 160268 307720 160274
rect 307668 160210 307720 160216
rect 307484 160132 307536 160138
rect 307484 160074 307536 160080
rect 307574 160032 307630 160041
rect 307574 159967 307630 159976
rect 307392 159384 307444 159390
rect 307392 159326 307444 159332
rect 307206 159080 307262 159089
rect 307206 159015 307262 159024
rect 307220 148374 307248 159015
rect 307588 158778 307616 159967
rect 307666 159624 307722 159633
rect 307666 159559 307722 159568
rect 307680 158846 307708 159559
rect 307668 158840 307720 158846
rect 307668 158782 307720 158788
rect 307576 158772 307628 158778
rect 307576 158714 307628 158720
rect 307666 158264 307722 158273
rect 307666 158199 307722 158208
rect 307298 157856 307354 157865
rect 307298 157791 307354 157800
rect 307312 157418 307340 157791
rect 307680 157554 307708 158199
rect 307668 157548 307720 157554
rect 307668 157490 307720 157496
rect 307666 157448 307722 157457
rect 307300 157412 307352 157418
rect 307666 157383 307722 157392
rect 307300 157354 307352 157360
rect 307680 156670 307708 157383
rect 307668 156664 307720 156670
rect 307482 156632 307538 156641
rect 307668 156606 307720 156612
rect 307482 156567 307538 156576
rect 307390 156224 307446 156233
rect 307390 156159 307446 156168
rect 307404 153882 307432 156159
rect 307496 156058 307524 156567
rect 307484 156052 307536 156058
rect 307484 155994 307536 156000
rect 307482 155680 307538 155689
rect 307482 155615 307538 155624
rect 307496 154630 307524 155615
rect 307574 155272 307630 155281
rect 307574 155207 307630 155216
rect 307588 154766 307616 155207
rect 307666 154864 307722 154873
rect 307666 154799 307722 154808
rect 307576 154760 307628 154766
rect 307576 154702 307628 154708
rect 307680 154698 307708 154799
rect 307668 154692 307720 154698
rect 307668 154634 307720 154640
rect 307484 154624 307536 154630
rect 307484 154566 307536 154572
rect 307482 154456 307538 154465
rect 307482 154391 307538 154400
rect 307392 153876 307444 153882
rect 307392 153818 307444 153824
rect 307496 153270 307524 154391
rect 307666 154048 307722 154057
rect 307666 153983 307722 153992
rect 307574 153640 307630 153649
rect 307574 153575 307630 153584
rect 307484 153264 307536 153270
rect 307484 153206 307536 153212
rect 307482 152688 307538 152697
rect 307482 152623 307538 152632
rect 307496 151910 307524 152623
rect 307588 152522 307616 153575
rect 307680 153338 307708 153983
rect 307668 153332 307720 153338
rect 307668 153274 307720 153280
rect 307576 152516 307628 152522
rect 307576 152458 307628 152464
rect 307484 151904 307536 151910
rect 307484 151846 307536 151852
rect 307666 151872 307722 151881
rect 307666 151807 307668 151816
rect 307720 151807 307722 151816
rect 307668 151778 307720 151784
rect 307482 151464 307538 151473
rect 307482 151399 307538 151408
rect 307390 150648 307446 150657
rect 307390 150583 307446 150592
rect 307298 149288 307354 149297
rect 307298 149223 307300 149232
rect 307352 149223 307354 149232
rect 307300 149194 307352 149200
rect 307208 148368 307260 148374
rect 307208 148310 307260 148316
rect 307114 148064 307170 148073
rect 307114 147999 307170 148008
rect 307024 145580 307076 145586
rect 307024 145522 307076 145528
rect 306930 144664 306986 144673
rect 306930 144599 306986 144608
rect 306562 144256 306618 144265
rect 306562 144191 306618 144200
rect 306576 141438 306604 144191
rect 306944 143614 306972 144599
rect 306932 143608 306984 143614
rect 306932 143550 306984 143556
rect 306746 143032 306802 143041
rect 306746 142967 306802 142976
rect 306760 142254 306788 142967
rect 306748 142248 306800 142254
rect 306748 142190 306800 142196
rect 306564 141432 306616 141438
rect 306564 141374 306616 141380
rect 307022 141264 307078 141273
rect 307022 141199 307078 141208
rect 306930 136640 306986 136649
rect 306930 136575 306986 136584
rect 306944 135318 306972 136575
rect 306932 135312 306984 135318
rect 306932 135254 306984 135260
rect 305734 134464 305790 134473
rect 305734 134399 305790 134408
rect 305644 126268 305696 126274
rect 305644 126210 305696 126216
rect 305642 124672 305698 124681
rect 305642 124607 305698 124616
rect 304540 120284 304592 120290
rect 304540 120226 304592 120232
rect 304354 115152 304410 115161
rect 304354 115087 304410 115096
rect 304448 114708 304500 114714
rect 304448 114650 304500 114656
rect 304264 110628 304316 110634
rect 304264 110570 304316 110576
rect 303160 108996 303212 109002
rect 303160 108938 303212 108944
rect 303068 107704 303120 107710
rect 303068 107646 303120 107652
rect 303080 60042 303108 107646
rect 303160 103692 303212 103698
rect 303160 103634 303212 103640
rect 303172 68338 303200 103634
rect 303160 68332 303212 68338
rect 303160 68274 303212 68280
rect 303068 60036 303120 60042
rect 303068 59978 303120 59984
rect 304276 40798 304304 110570
rect 304356 109200 304408 109206
rect 304356 109142 304408 109148
rect 304368 53174 304396 109142
rect 304460 71058 304488 114650
rect 304552 76566 304580 120226
rect 304540 76560 304592 76566
rect 304540 76502 304592 76508
rect 304448 71052 304500 71058
rect 304448 70994 304500 71000
rect 304356 53168 304408 53174
rect 304356 53110 304408 53116
rect 304264 40792 304316 40798
rect 304264 40734 304316 40740
rect 302976 24200 303028 24206
rect 302976 24142 303028 24148
rect 302884 17332 302936 17338
rect 302884 17274 302936 17280
rect 305656 15910 305684 124607
rect 305748 73914 305776 134399
rect 306930 133648 306986 133657
rect 306930 133583 306986 133592
rect 306562 133240 306618 133249
rect 306562 133175 306618 133184
rect 306576 132530 306604 133175
rect 306944 132598 306972 133583
rect 306932 132592 306984 132598
rect 306932 132534 306984 132540
rect 306564 132524 306616 132530
rect 306564 132466 306616 132472
rect 306930 132288 306986 132297
rect 306930 132223 306986 132232
rect 306944 131170 306972 132223
rect 306932 131164 306984 131170
rect 306932 131106 306984 131112
rect 306746 129296 306802 129305
rect 306746 129231 306802 129240
rect 306760 128382 306788 129231
rect 306748 128376 306800 128382
rect 306748 128318 306800 128324
rect 306562 126440 306618 126449
rect 306562 126375 306618 126384
rect 306576 125730 306604 126375
rect 306930 125896 306986 125905
rect 306930 125831 306986 125840
rect 306564 125724 306616 125730
rect 306564 125666 306616 125672
rect 306944 125662 306972 125831
rect 306932 125656 306984 125662
rect 306932 125598 306984 125604
rect 306930 125488 306986 125497
rect 306930 125423 306986 125432
rect 306944 124438 306972 125423
rect 306932 124432 306984 124438
rect 306932 124374 306984 124380
rect 306930 121680 306986 121689
rect 306930 121615 306986 121624
rect 306944 121514 306972 121615
rect 306932 121508 306984 121514
rect 306932 121450 306984 121456
rect 306746 121272 306802 121281
rect 306746 121207 306802 121216
rect 306760 120222 306788 121207
rect 306748 120216 306800 120222
rect 306748 120158 306800 120164
rect 306930 120048 306986 120057
rect 306930 119983 306986 119992
rect 306562 119640 306618 119649
rect 306562 119575 306618 119584
rect 306576 118862 306604 119575
rect 306564 118856 306616 118862
rect 306564 118798 306616 118804
rect 306944 118726 306972 119983
rect 307036 119406 307064 141199
rect 307128 133210 307156 147999
rect 307298 147656 307354 147665
rect 307298 147591 307354 147600
rect 307206 145480 307262 145489
rect 307206 145415 307262 145424
rect 307116 133204 307168 133210
rect 307116 133146 307168 133152
rect 307114 130656 307170 130665
rect 307114 130591 307170 130600
rect 307024 119400 307076 119406
rect 307024 119342 307076 119348
rect 306932 118720 306984 118726
rect 306932 118662 306984 118668
rect 306562 118280 306618 118289
rect 306562 118215 306618 118224
rect 306576 117366 306604 118215
rect 306564 117360 306616 117366
rect 306564 117302 306616 117308
rect 306746 117056 306802 117065
rect 306746 116991 306802 117000
rect 306760 116074 306788 116991
rect 306748 116068 306800 116074
rect 306748 116010 306800 116016
rect 306746 115696 306802 115705
rect 306746 115631 306802 115640
rect 306760 114714 306788 115631
rect 306748 114708 306800 114714
rect 306748 114650 306800 114656
rect 307022 114064 307078 114073
rect 307022 113999 307078 114008
rect 306930 108080 306986 108089
rect 306930 108015 306986 108024
rect 305826 107808 305882 107817
rect 305826 107743 305882 107752
rect 305736 73908 305788 73914
rect 305736 73850 305788 73856
rect 305840 57254 305868 107743
rect 306944 107710 306972 108015
rect 306932 107704 306984 107710
rect 306932 107646 306984 107652
rect 305918 105224 305974 105233
rect 305918 105159 305974 105168
rect 305932 65550 305960 105159
rect 306746 103456 306802 103465
rect 306746 103391 306802 103400
rect 306760 102338 306788 103391
rect 306748 102332 306800 102338
rect 306748 102274 306800 102280
rect 306562 101688 306618 101697
rect 306562 101623 306618 101632
rect 306576 100842 306604 101623
rect 306564 100836 306616 100842
rect 306564 100778 306616 100784
rect 306746 97880 306802 97889
rect 306746 97815 306802 97824
rect 306760 96830 306788 97815
rect 306748 96824 306800 96830
rect 306748 96766 306800 96772
rect 305920 65544 305972 65550
rect 305920 65486 305972 65492
rect 305828 57248 305880 57254
rect 305828 57190 305880 57196
rect 307036 28286 307064 113999
rect 307128 47598 307156 130591
rect 307220 127634 307248 145415
rect 307312 144226 307340 147591
rect 307300 144220 307352 144226
rect 307300 144162 307352 144168
rect 307298 142488 307354 142497
rect 307298 142423 307354 142432
rect 307312 134570 307340 142423
rect 307404 142322 307432 150583
rect 307496 150550 307524 151399
rect 307666 151056 307722 151065
rect 307666 150991 307722 151000
rect 307484 150544 307536 150550
rect 307484 150486 307536 150492
rect 307680 150482 307708 150991
rect 307668 150476 307720 150482
rect 307668 150418 307720 150424
rect 307482 149832 307538 149841
rect 307482 149767 307538 149776
rect 307496 149122 307524 149767
rect 307484 149116 307536 149122
rect 307484 149058 307536 149064
rect 307666 148880 307722 148889
rect 307666 148815 307722 148824
rect 307482 148472 307538 148481
rect 307482 148407 307538 148416
rect 307496 147762 307524 148407
rect 307484 147756 307536 147762
rect 307484 147698 307536 147704
rect 307680 147694 307708 148815
rect 307668 147688 307720 147694
rect 307668 147630 307720 147636
rect 307666 146840 307722 146849
rect 307666 146775 307722 146784
rect 307680 146470 307708 146775
rect 307668 146464 307720 146470
rect 307574 146432 307630 146441
rect 307668 146406 307720 146412
rect 307574 146367 307630 146376
rect 307588 146334 307616 146367
rect 307576 146328 307628 146334
rect 307576 146270 307628 146276
rect 307482 145888 307538 145897
rect 307482 145823 307538 145832
rect 307496 145042 307524 145823
rect 307666 145072 307722 145081
rect 307484 145036 307536 145042
rect 307666 145007 307722 145016
rect 307484 144978 307536 144984
rect 307680 144974 307708 145007
rect 307668 144968 307720 144974
rect 307668 144910 307720 144916
rect 307482 143848 307538 143857
rect 307482 143783 307538 143792
rect 307496 143682 307524 143783
rect 307484 143676 307536 143682
rect 307484 143618 307536 143624
rect 307666 143440 307722 143449
rect 307666 143375 307722 143384
rect 307392 142316 307444 142322
rect 307392 142258 307444 142264
rect 307680 142186 307708 143375
rect 307668 142180 307720 142186
rect 307668 142122 307720 142128
rect 307574 142080 307630 142089
rect 307574 142015 307630 142024
rect 307482 141672 307538 141681
rect 307482 141607 307538 141616
rect 307496 140826 307524 141607
rect 307588 140894 307616 142015
rect 307668 140956 307720 140962
rect 307668 140898 307720 140904
rect 307576 140888 307628 140894
rect 307680 140865 307708 140898
rect 307576 140830 307628 140836
rect 307666 140856 307722 140865
rect 307484 140820 307536 140826
rect 307666 140791 307722 140800
rect 307484 140762 307536 140768
rect 307666 139632 307722 139641
rect 307666 139567 307722 139576
rect 307680 139466 307708 139567
rect 307668 139460 307720 139466
rect 307668 139402 307720 139408
rect 307482 139088 307538 139097
rect 307482 139023 307538 139032
rect 307496 138038 307524 139023
rect 307574 138680 307630 138689
rect 307574 138615 307630 138624
rect 307588 138106 307616 138615
rect 307666 138272 307722 138281
rect 307666 138207 307722 138216
rect 307680 138174 307708 138207
rect 307668 138168 307720 138174
rect 307668 138110 307720 138116
rect 307576 138100 307628 138106
rect 307576 138042 307628 138048
rect 307484 138032 307536 138038
rect 307484 137974 307536 137980
rect 307574 137864 307630 137873
rect 307574 137799 307630 137808
rect 307482 137456 307538 137465
rect 307482 137391 307538 137400
rect 307496 136814 307524 137391
rect 307484 136808 307536 136814
rect 307484 136750 307536 136756
rect 307588 136746 307616 137799
rect 307666 137048 307722 137057
rect 307666 136983 307722 136992
rect 307576 136740 307628 136746
rect 307576 136682 307628 136688
rect 307680 136678 307708 136983
rect 307668 136672 307720 136678
rect 307668 136614 307720 136620
rect 307482 136232 307538 136241
rect 307482 136167 307538 136176
rect 307496 135454 307524 136167
rect 307666 135688 307722 135697
rect 307666 135623 307722 135632
rect 307484 135448 307536 135454
rect 307484 135390 307536 135396
rect 307680 135386 307708 135623
rect 307668 135380 307720 135386
rect 307668 135322 307720 135328
rect 307482 134872 307538 134881
rect 307482 134807 307538 134816
rect 307300 134564 307352 134570
rect 307300 134506 307352 134512
rect 307496 134094 307524 134807
rect 307484 134088 307536 134094
rect 307484 134030 307536 134036
rect 307666 134056 307722 134065
rect 307666 133991 307668 134000
rect 307720 133991 307722 134000
rect 307668 133962 307720 133968
rect 307666 132696 307722 132705
rect 307666 132631 307668 132640
rect 307720 132631 307722 132640
rect 307668 132602 307720 132608
rect 307666 131880 307722 131889
rect 307666 131815 307722 131824
rect 307390 131472 307446 131481
rect 307390 131407 307446 131416
rect 307300 129872 307352 129878
rect 307298 129840 307300 129849
rect 307352 129840 307354 129849
rect 307298 129775 307354 129784
rect 307298 128480 307354 128489
rect 307298 128415 307300 128424
rect 307352 128415 307354 128424
rect 307300 128386 307352 128392
rect 307208 127628 307260 127634
rect 307208 127570 307260 127576
rect 307404 122834 307432 131407
rect 307680 131238 307708 131815
rect 307668 131232 307720 131238
rect 307668 131174 307720 131180
rect 307666 130248 307722 130257
rect 307666 130183 307722 130192
rect 307680 129810 307708 130183
rect 307668 129804 307720 129810
rect 307668 129746 307720 129752
rect 307666 128888 307722 128897
rect 307666 128823 307722 128832
rect 307680 128518 307708 128823
rect 307668 128512 307720 128518
rect 307668 128454 307720 128460
rect 307574 127664 307630 127673
rect 307574 127599 307630 127608
rect 307588 127090 307616 127599
rect 307666 127256 307722 127265
rect 307666 127191 307722 127200
rect 307576 127084 307628 127090
rect 307576 127026 307628 127032
rect 307680 127022 307708 127191
rect 307668 127016 307720 127022
rect 307668 126958 307720 126964
rect 307482 125080 307538 125089
rect 307482 125015 307538 125024
rect 307496 124234 307524 125015
rect 307668 124296 307720 124302
rect 307666 124264 307668 124273
rect 307720 124264 307722 124273
rect 307484 124228 307536 124234
rect 307666 124199 307722 124208
rect 307484 124170 307536 124176
rect 307574 123856 307630 123865
rect 307574 123791 307630 123800
rect 307482 123040 307538 123049
rect 307588 123010 307616 123791
rect 307666 123448 307722 123457
rect 307666 123383 307722 123392
rect 307482 122975 307538 122984
rect 307576 123004 307628 123010
rect 307496 122874 307524 122975
rect 307576 122946 307628 122952
rect 307680 122942 307708 123383
rect 307668 122936 307720 122942
rect 307668 122878 307720 122884
rect 307312 122806 307432 122834
rect 307484 122868 307536 122874
rect 307484 122810 307536 122816
rect 307206 96248 307262 96257
rect 307206 96183 307262 96192
rect 307220 51746 307248 96183
rect 307312 87650 307340 122806
rect 307482 122496 307538 122505
rect 307482 122431 307538 122440
rect 307496 121650 307524 122431
rect 307666 122088 307722 122097
rect 307666 122023 307722 122032
rect 307484 121644 307536 121650
rect 307484 121586 307536 121592
rect 307680 121582 307708 122023
rect 307668 121576 307720 121582
rect 307668 121518 307720 121524
rect 307482 120864 307538 120873
rect 307482 120799 307538 120808
rect 307496 120290 307524 120799
rect 307666 120456 307722 120465
rect 307666 120391 307722 120400
rect 307484 120284 307536 120290
rect 307484 120226 307536 120232
rect 307680 120154 307708 120391
rect 307668 120148 307720 120154
rect 307668 120090 307720 120096
rect 307666 119096 307722 119105
rect 307666 119031 307722 119040
rect 307680 118794 307708 119031
rect 307668 118788 307720 118794
rect 307668 118730 307720 118736
rect 307574 118688 307630 118697
rect 307574 118623 307630 118632
rect 307588 117502 307616 118623
rect 307666 117872 307722 117881
rect 307666 117807 307722 117816
rect 307576 117496 307628 117502
rect 307576 117438 307628 117444
rect 307680 117434 307708 117807
rect 307668 117428 307720 117434
rect 307668 117370 307720 117376
rect 307574 116648 307630 116657
rect 307574 116583 307630 116592
rect 307588 116006 307616 116583
rect 307666 116240 307722 116249
rect 307666 116175 307722 116184
rect 307680 116142 307708 116175
rect 307668 116136 307720 116142
rect 307668 116078 307720 116084
rect 307576 116000 307628 116006
rect 307576 115942 307628 115948
rect 307574 115288 307630 115297
rect 307574 115223 307630 115232
rect 307588 114646 307616 115223
rect 307666 114880 307722 114889
rect 307666 114815 307722 114824
rect 307576 114640 307628 114646
rect 307576 114582 307628 114588
rect 307680 114578 307708 114815
rect 307668 114572 307720 114578
rect 307668 114514 307720 114520
rect 307574 113656 307630 113665
rect 307574 113591 307630 113600
rect 307588 113218 307616 113591
rect 307668 113280 307720 113286
rect 307666 113248 307668 113257
rect 307720 113248 307722 113257
rect 307576 113212 307628 113218
rect 307666 113183 307722 113192
rect 307576 113154 307628 113160
rect 307482 112704 307538 112713
rect 307482 112639 307538 112648
rect 307496 111926 307524 112639
rect 307574 112296 307630 112305
rect 307574 112231 307630 112240
rect 307484 111920 307536 111926
rect 307484 111862 307536 111868
rect 307588 111858 307616 112231
rect 307668 111988 307720 111994
rect 307668 111930 307720 111936
rect 307680 111897 307708 111930
rect 307666 111888 307722 111897
rect 307576 111852 307628 111858
rect 307666 111823 307722 111832
rect 307576 111794 307628 111800
rect 307482 111480 307538 111489
rect 307482 111415 307538 111424
rect 307496 110566 307524 111415
rect 307666 111072 307722 111081
rect 307666 111007 307722 111016
rect 307574 110664 307630 110673
rect 307680 110634 307708 111007
rect 307574 110599 307630 110608
rect 307668 110628 307720 110634
rect 307484 110560 307536 110566
rect 307484 110502 307536 110508
rect 307588 110498 307616 110599
rect 307668 110570 307720 110576
rect 307576 110492 307628 110498
rect 307576 110434 307628 110440
rect 307482 110256 307538 110265
rect 307482 110191 307538 110200
rect 307496 109206 307524 110191
rect 307574 109848 307630 109857
rect 307574 109783 307630 109792
rect 307484 109200 307536 109206
rect 307484 109142 307536 109148
rect 307588 109138 307616 109783
rect 307666 109304 307722 109313
rect 307666 109239 307722 109248
rect 307576 109132 307628 109138
rect 307576 109074 307628 109080
rect 307680 109070 307708 109239
rect 307668 109064 307720 109070
rect 307668 109006 307720 109012
rect 307482 108896 307538 108905
rect 307482 108831 307538 108840
rect 307496 107817 307524 108831
rect 307574 108488 307630 108497
rect 307574 108423 307630 108432
rect 307482 107808 307538 107817
rect 307588 107778 307616 108423
rect 307668 107908 307720 107914
rect 307668 107850 307720 107856
rect 307482 107743 307538 107752
rect 307576 107772 307628 107778
rect 307576 107714 307628 107720
rect 307680 107681 307708 107850
rect 307666 107672 307722 107681
rect 307666 107607 307722 107616
rect 307482 107264 307538 107273
rect 307482 107199 307538 107208
rect 307496 106486 307524 107199
rect 307574 106856 307630 106865
rect 307574 106791 307630 106800
rect 307484 106480 307536 106486
rect 307484 106422 307536 106428
rect 307588 106418 307616 106791
rect 307666 106448 307722 106457
rect 307576 106412 307628 106418
rect 307666 106383 307722 106392
rect 307576 106354 307628 106360
rect 307680 106350 307708 106383
rect 307668 106344 307720 106350
rect 307668 106286 307720 106292
rect 307666 105904 307722 105913
rect 307666 105839 307722 105848
rect 307482 105496 307538 105505
rect 307482 105431 307538 105440
rect 307496 105058 307524 105431
rect 307680 105233 307708 105839
rect 307666 105224 307722 105233
rect 307666 105159 307722 105168
rect 307666 105088 307722 105097
rect 307484 105052 307536 105058
rect 307666 105023 307722 105032
rect 307484 104994 307536 105000
rect 307680 104990 307708 105023
rect 307668 104984 307720 104990
rect 307668 104926 307720 104932
rect 307574 104680 307630 104689
rect 307574 104615 307630 104624
rect 307482 104272 307538 104281
rect 307482 104207 307538 104216
rect 307496 103562 307524 104207
rect 307588 103698 307616 104615
rect 307666 103864 307722 103873
rect 307666 103799 307722 103808
rect 307576 103692 307628 103698
rect 307576 103634 307628 103640
rect 307680 103630 307708 103799
rect 307668 103624 307720 103630
rect 307668 103566 307720 103572
rect 307484 103556 307536 103562
rect 307484 103498 307536 103504
rect 307482 103048 307538 103057
rect 307482 102983 307538 102992
rect 307496 102202 307524 102983
rect 307666 102504 307722 102513
rect 307666 102439 307722 102448
rect 307680 102270 307708 102439
rect 307668 102264 307720 102270
rect 307668 102206 307720 102212
rect 307484 102196 307536 102202
rect 307484 102138 307536 102144
rect 308218 102096 308274 102105
rect 308218 102031 308274 102040
rect 308232 101153 308260 102031
rect 308218 101144 308274 101153
rect 308218 101079 308274 101088
rect 307666 100872 307722 100881
rect 307666 100807 307722 100816
rect 307680 100774 307708 100807
rect 307668 100768 307720 100774
rect 307668 100710 307720 100716
rect 307574 100464 307630 100473
rect 307574 100399 307630 100408
rect 307588 99482 307616 100399
rect 307666 99648 307722 99657
rect 307666 99583 307722 99592
rect 307576 99476 307628 99482
rect 307576 99418 307628 99424
rect 307680 99414 307708 99583
rect 307668 99408 307720 99414
rect 307668 99350 307720 99356
rect 307666 99104 307722 99113
rect 307666 99039 307722 99048
rect 307574 98696 307630 98705
rect 307574 98631 307630 98640
rect 307482 98288 307538 98297
rect 307482 98223 307538 98232
rect 307496 98122 307524 98223
rect 307484 98116 307536 98122
rect 307484 98058 307536 98064
rect 307588 98054 307616 98631
rect 307680 98190 307708 99039
rect 307668 98184 307720 98190
rect 307668 98126 307720 98132
rect 307576 98048 307628 98054
rect 307576 97990 307628 97996
rect 307482 97472 307538 97481
rect 307482 97407 307538 97416
rect 307496 96694 307524 97407
rect 307668 96756 307720 96762
rect 307668 96698 307720 96704
rect 307484 96688 307536 96694
rect 307680 96665 307708 96698
rect 307484 96630 307536 96636
rect 307666 96656 307722 96665
rect 307666 96591 307722 96600
rect 307300 87644 307352 87650
rect 307300 87586 307352 87592
rect 308416 76566 308444 357750
rect 308588 285728 308640 285734
rect 308588 285670 308640 285676
rect 308496 207868 308548 207874
rect 308496 207810 308548 207816
rect 308404 76560 308456 76566
rect 308404 76502 308456 76508
rect 307208 51740 307260 51746
rect 307208 51682 307260 51688
rect 307116 47592 307168 47598
rect 307116 47534 307168 47540
rect 307024 28280 307076 28286
rect 307024 28222 307076 28228
rect 305644 15904 305696 15910
rect 305644 15846 305696 15852
rect 306380 14612 306432 14618
rect 306380 14554 306432 14560
rect 301962 6216 302018 6225
rect 301504 6180 301556 6186
rect 301962 6151 302018 6160
rect 305552 6180 305604 6186
rect 301504 6122 301556 6128
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 300780 480 300808 3470
rect 301976 480 302004 6151
rect 305552 6122 305604 6128
rect 304356 4888 304408 4894
rect 304356 4830 304408 4836
rect 303158 3496 303214 3505
rect 303158 3431 303214 3440
rect 303172 480 303200 3431
rect 304368 480 304396 4830
rect 305564 480 305592 6122
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 354 306420 14554
rect 307942 3496 307998 3505
rect 307942 3431 307998 3440
rect 307956 480 307984 3431
rect 308508 3194 308536 207810
rect 308600 90370 308628 285670
rect 309152 240038 309180 402222
rect 310520 362976 310572 362982
rect 310520 362918 310572 362924
rect 309784 360460 309836 360466
rect 309784 360402 309836 360408
rect 309692 260908 309744 260914
rect 309692 260850 309744 260856
rect 309140 240032 309192 240038
rect 309140 239974 309192 239980
rect 308678 140040 308734 140049
rect 308678 139975 308734 139984
rect 308692 139505 308720 139975
rect 308678 139496 308734 139505
rect 308678 139431 308734 139440
rect 309704 90438 309732 260850
rect 309692 90432 309744 90438
rect 309692 90374 309744 90380
rect 308588 90364 308640 90370
rect 308588 90306 308640 90312
rect 309046 4040 309102 4049
rect 309046 3975 309102 3984
rect 308496 3188 308548 3194
rect 308496 3130 308548 3136
rect 309060 480 309088 3975
rect 309796 3466 309824 360402
rect 309876 339516 309928 339522
rect 309876 339458 309928 339464
rect 309888 73710 309916 339458
rect 310428 240032 310480 240038
rect 310428 239974 310480 239980
rect 310440 239426 310468 239974
rect 310428 239420 310480 239426
rect 310428 239362 310480 239368
rect 310532 177410 310560 362918
rect 310624 238678 310652 408478
rect 312544 360392 312596 360398
rect 312544 360334 312596 360340
rect 311164 253972 311216 253978
rect 311164 253914 311216 253920
rect 310612 238672 310664 238678
rect 310612 238614 310664 238620
rect 311176 232626 311204 253914
rect 311164 232620 311216 232626
rect 311164 232562 311216 232568
rect 311164 218748 311216 218754
rect 311164 218690 311216 218696
rect 311176 177478 311204 218690
rect 311256 198076 311308 198082
rect 311256 198018 311308 198024
rect 311268 178770 311296 198018
rect 311256 178764 311308 178770
rect 311256 178706 311308 178712
rect 312556 178702 312584 360334
rect 313292 238610 313320 536046
rect 313372 357740 313424 357746
rect 313372 357682 313424 357688
rect 313280 238604 313332 238610
rect 313280 238546 313332 238552
rect 313384 232558 313412 357682
rect 314672 238785 314700 556174
rect 328460 539640 328512 539646
rect 328460 539582 328512 539588
rect 324964 502376 325016 502382
rect 324964 502318 325016 502324
rect 317420 474768 317472 474774
rect 317420 474710 317472 474716
rect 315304 393372 315356 393378
rect 315304 393314 315356 393320
rect 314658 238776 314714 238785
rect 314658 238711 314714 238720
rect 314566 235240 314622 235249
rect 314566 235175 314622 235184
rect 313372 232552 313424 232558
rect 313372 232494 313424 232500
rect 313924 211812 313976 211818
rect 313924 211754 313976 211760
rect 313832 181484 313884 181490
rect 313832 181426 313884 181432
rect 312544 178696 312596 178702
rect 312544 178638 312596 178644
rect 311164 177472 311216 177478
rect 311164 177414 311216 177420
rect 310520 177404 310572 177410
rect 310520 177346 310572 177352
rect 313844 176662 313872 181426
rect 313936 177410 313964 211754
rect 314580 181490 314608 235175
rect 314568 181484 314620 181490
rect 314568 181426 314620 181432
rect 315316 180130 315344 393314
rect 317432 234530 317460 474710
rect 322940 420980 322992 420986
rect 322940 420922 322992 420928
rect 319444 395344 319496 395350
rect 319444 395286 319496 395292
rect 317420 234524 317472 234530
rect 317420 234466 317472 234472
rect 318064 234524 318116 234530
rect 318064 234466 318116 234472
rect 315396 217320 315448 217326
rect 315396 217262 315448 217268
rect 315304 180124 315356 180130
rect 315304 180066 315356 180072
rect 313924 177404 313976 177410
rect 313924 177346 313976 177352
rect 313832 176656 313884 176662
rect 313832 176598 313884 176604
rect 315408 175982 315436 217262
rect 315488 191140 315540 191146
rect 315488 191082 315540 191088
rect 315500 177546 315528 191082
rect 318076 181694 318104 234466
rect 318156 207664 318208 207670
rect 318156 207606 318208 207612
rect 318064 181688 318116 181694
rect 318064 181630 318116 181636
rect 316040 178084 316092 178090
rect 316040 178026 316092 178032
rect 315488 177540 315540 177546
rect 315488 177482 315540 177488
rect 315396 175976 315448 175982
rect 316052 175930 316080 178026
rect 318168 177449 318196 207606
rect 318248 200864 318300 200870
rect 318248 200806 318300 200812
rect 318154 177440 318210 177449
rect 318154 177375 318210 177384
rect 318260 176225 318288 200806
rect 318432 185700 318484 185706
rect 318432 185642 318484 185648
rect 318444 176633 318472 185642
rect 319456 184414 319484 395286
rect 322952 237386 322980 420922
rect 323032 385688 323084 385694
rect 323032 385630 323084 385636
rect 322940 237380 322992 237386
rect 322940 237322 322992 237328
rect 322952 236026 322980 237322
rect 322940 236020 322992 236026
rect 322940 235962 322992 235968
rect 323044 235249 323072 385630
rect 323584 236020 323636 236026
rect 323584 235962 323636 235968
rect 323030 235240 323086 235249
rect 323030 235175 323086 235184
rect 322940 213240 322992 213246
rect 322940 213182 322992 213188
rect 321652 209160 321704 209166
rect 321652 209102 321704 209108
rect 321560 192568 321612 192574
rect 321560 192510 321612 192516
rect 319536 188352 319588 188358
rect 319536 188294 319588 188300
rect 319444 184408 319496 184414
rect 319444 184350 319496 184356
rect 318430 176624 318486 176633
rect 319548 176594 319576 188294
rect 321284 185632 321336 185638
rect 321284 185574 321336 185580
rect 318430 176559 318486 176568
rect 319536 176588 319588 176594
rect 319536 176530 319588 176536
rect 318246 176216 318302 176225
rect 318246 176151 318302 176160
rect 315396 175918 315448 175924
rect 316020 175902 316080 175930
rect 321296 170377 321324 185574
rect 321468 176656 321520 176662
rect 321468 176598 321520 176604
rect 321480 176089 321508 176598
rect 321466 176080 321522 176089
rect 321466 176015 321522 176024
rect 321282 170368 321338 170377
rect 321282 170303 321338 170312
rect 321572 106049 321600 192510
rect 321664 148345 321692 209102
rect 321836 186992 321888 186998
rect 321836 186934 321888 186940
rect 321744 176588 321796 176594
rect 321744 176530 321796 176536
rect 321756 174457 321784 176530
rect 321742 174448 321798 174457
rect 321742 174383 321798 174392
rect 321848 172689 321876 186934
rect 321834 172680 321890 172689
rect 321834 172615 321890 172624
rect 321650 148336 321706 148345
rect 321650 148271 321706 148280
rect 321650 107536 321706 107545
rect 321650 107471 321706 107480
rect 321558 106040 321614 106049
rect 321558 105975 321614 105984
rect 321558 102232 321614 102241
rect 321558 102167 321614 102176
rect 321374 97336 321430 97345
rect 321374 97271 321430 97280
rect 321388 95985 321416 97271
rect 321374 95976 321430 95985
rect 321374 95911 321430 95920
rect 321466 95840 321522 95849
rect 318064 95804 318116 95810
rect 321466 95775 321468 95784
rect 318064 95746 318116 95752
rect 321520 95775 321522 95784
rect 321468 95746 321520 95752
rect 313280 83496 313332 83502
rect 313280 83438 313332 83444
rect 310518 79384 310574 79393
rect 310518 79319 310574 79328
rect 309876 73704 309928 73710
rect 309876 73646 309928 73652
rect 310532 16574 310560 79319
rect 311900 31204 311952 31210
rect 311900 31146 311952 31152
rect 311912 16574 311940 31146
rect 313292 16574 313320 83438
rect 318076 78674 318104 95746
rect 321572 93770 321600 102167
rect 321664 95130 321692 107471
rect 322952 106321 322980 213182
rect 323030 176624 323086 176633
rect 323030 176559 323086 176568
rect 323044 173233 323072 176559
rect 323030 173224 323086 173233
rect 323030 173159 323086 173168
rect 323596 137358 323624 235962
rect 324596 233912 324648 233918
rect 324596 233854 324648 233860
rect 324318 223680 324374 223689
rect 324318 223615 324374 223624
rect 324332 223582 324360 223615
rect 324320 223576 324372 223582
rect 324320 223518 324372 223524
rect 324410 193896 324466 193905
rect 324410 193831 324466 193840
rect 323676 186992 323728 186998
rect 323676 186934 323728 186940
rect 323688 146305 323716 186934
rect 324320 170944 324372 170950
rect 324318 170912 324320 170921
rect 324372 170912 324374 170921
rect 324318 170847 324374 170856
rect 324320 169720 324372 169726
rect 324320 169662 324372 169668
rect 324332 168609 324360 169662
rect 324318 168600 324374 168609
rect 324318 168535 324374 168544
rect 324320 168360 324372 168366
rect 324320 168302 324372 168308
rect 324332 167113 324360 168302
rect 324424 167793 324452 193831
rect 324504 187128 324556 187134
rect 324504 187070 324556 187076
rect 324516 174729 324544 187070
rect 324502 174720 324558 174729
rect 324502 174655 324558 174664
rect 324410 167784 324466 167793
rect 324410 167719 324466 167728
rect 324318 167104 324374 167113
rect 324318 167039 324374 167048
rect 324412 165572 324464 165578
rect 324412 165514 324464 165520
rect 324320 165504 324372 165510
rect 324318 165472 324320 165481
rect 324372 165472 324374 165481
rect 324318 165407 324374 165416
rect 324424 164801 324452 165514
rect 324410 164792 324466 164801
rect 324410 164727 324466 164736
rect 324320 164212 324372 164218
rect 324320 164154 324372 164160
rect 324332 163985 324360 164154
rect 324412 164144 324464 164150
rect 324412 164086 324464 164092
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324424 163169 324452 164086
rect 324410 163160 324466 163169
rect 324410 163095 324466 163104
rect 324320 162852 324372 162858
rect 324320 162794 324372 162800
rect 324332 161673 324360 162794
rect 324318 161664 324374 161673
rect 324318 161599 324374 161608
rect 324320 161424 324372 161430
rect 324320 161366 324372 161372
rect 324332 160177 324360 161366
rect 324318 160168 324374 160177
rect 324318 160103 324374 160112
rect 324320 160064 324372 160070
rect 324320 160006 324372 160012
rect 324332 159361 324360 160006
rect 324318 159352 324374 159361
rect 324318 159287 324374 159296
rect 324412 158704 324464 158710
rect 324412 158646 324464 158652
rect 324320 158636 324372 158642
rect 324320 158578 324372 158584
rect 324332 158545 324360 158578
rect 324318 158536 324374 158545
rect 324318 158471 324374 158480
rect 324424 157865 324452 158646
rect 324410 157856 324466 157865
rect 324410 157791 324466 157800
rect 324320 157344 324372 157350
rect 324320 157286 324372 157292
rect 324332 157049 324360 157286
rect 324412 157208 324464 157214
rect 324412 157150 324464 157156
rect 324318 157040 324374 157049
rect 324318 156975 324374 156984
rect 324424 156369 324452 157150
rect 324410 156360 324466 156369
rect 324410 156295 324466 156304
rect 324320 155916 324372 155922
rect 324320 155858 324372 155864
rect 324332 154737 324360 155858
rect 324608 155553 324636 233854
rect 324976 223689 325004 502318
rect 327264 434784 327316 434790
rect 327264 434726 327316 434732
rect 325056 324352 325108 324358
rect 325056 324294 325108 324300
rect 325068 283626 325096 324294
rect 325056 283620 325108 283626
rect 325056 283562 325108 283568
rect 325056 264988 325108 264994
rect 325056 264930 325108 264936
rect 325068 225622 325096 264930
rect 325148 249824 325200 249830
rect 325148 249766 325200 249772
rect 325056 225616 325108 225622
rect 325056 225558 325108 225564
rect 324962 223680 325018 223689
rect 324962 223615 325018 223624
rect 325160 222902 325188 249766
rect 327172 238060 327224 238066
rect 327172 238002 327224 238008
rect 325792 231124 325844 231130
rect 325792 231066 325844 231072
rect 325148 222896 325200 222902
rect 325148 222838 325200 222844
rect 325698 210352 325754 210361
rect 325698 210287 325754 210296
rect 324594 155544 324650 155553
rect 324594 155479 324650 155488
rect 324318 154728 324374 154737
rect 324318 154663 324374 154672
rect 324320 154556 324372 154562
rect 324320 154498 324372 154504
rect 324332 154057 324360 154498
rect 324412 154488 324464 154494
rect 324412 154430 324464 154436
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 324424 153241 324452 154430
rect 324410 153232 324466 153241
rect 324320 153196 324372 153202
rect 324410 153167 324466 153176
rect 324320 153138 324372 153144
rect 324332 152425 324360 153138
rect 324318 152416 324374 152425
rect 324318 152351 324374 152360
rect 324412 151768 324464 151774
rect 324318 151736 324374 151745
rect 324412 151710 324464 151716
rect 324318 151671 324320 151680
rect 324372 151671 324374 151680
rect 324320 151642 324372 151648
rect 324424 150929 324452 151710
rect 324410 150920 324466 150929
rect 324410 150855 324466 150864
rect 324320 150408 324372 150414
rect 324320 150350 324372 150356
rect 324332 149433 324360 150350
rect 324318 149424 324374 149433
rect 324318 149359 324374 149368
rect 324320 149048 324372 149054
rect 324320 148990 324372 148996
rect 324332 148617 324360 148990
rect 324318 148608 324374 148617
rect 324318 148543 324374 148552
rect 324320 147620 324372 147626
rect 324320 147562 324372 147568
rect 324332 147121 324360 147562
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 323674 146296 323730 146305
rect 323674 146231 323730 146240
rect 324320 144900 324372 144906
rect 324320 144842 324372 144848
rect 324332 144809 324360 144842
rect 324318 144800 324374 144809
rect 324318 144735 324374 144744
rect 324320 143540 324372 143546
rect 324320 143482 324372 143488
rect 324332 143177 324360 143482
rect 324318 143168 324374 143177
rect 324318 143103 324374 143112
rect 324320 139392 324372 139398
rect 324320 139334 324372 139340
rect 324332 138553 324360 139334
rect 324318 138544 324374 138553
rect 324318 138479 324374 138488
rect 324320 137964 324372 137970
rect 324320 137906 324372 137912
rect 324332 137873 324360 137906
rect 324504 137896 324556 137902
rect 324318 137864 324374 137873
rect 324504 137838 324556 137844
rect 324318 137799 324374 137808
rect 323584 137352 323636 137358
rect 323584 137294 323636 137300
rect 324412 137352 324464 137358
rect 324412 137294 324464 137300
rect 324320 135244 324372 135250
rect 324320 135186 324372 135192
rect 324332 134745 324360 135186
rect 324318 134736 324374 134745
rect 324318 134671 324374 134680
rect 324320 133884 324372 133890
rect 324320 133826 324372 133832
rect 324332 133249 324360 133826
rect 324318 133240 324374 133249
rect 324318 133175 324374 133184
rect 324424 132494 324452 137294
rect 324516 137057 324544 137838
rect 324502 137048 324558 137057
rect 324502 136983 324558 136992
rect 324504 135176 324556 135182
rect 324504 135118 324556 135124
rect 324516 134065 324544 135118
rect 324502 134056 324558 134065
rect 324502 133991 324558 134000
rect 324424 132466 324544 132494
rect 324320 132456 324372 132462
rect 324318 132424 324320 132433
rect 324372 132424 324374 132433
rect 324318 132359 324374 132368
rect 324410 131744 324466 131753
rect 324410 131679 324466 131688
rect 324320 131096 324372 131102
rect 324320 131038 324372 131044
rect 324332 130121 324360 131038
rect 324424 130937 324452 131679
rect 324410 130928 324466 130937
rect 324410 130863 324466 130872
rect 324318 130112 324374 130121
rect 324318 130047 324374 130056
rect 324412 129736 324464 129742
rect 324412 129678 324464 129684
rect 324320 129668 324372 129674
rect 324320 129610 324372 129616
rect 324332 129441 324360 129610
rect 324318 129432 324374 129441
rect 324318 129367 324374 129376
rect 324424 128625 324452 129678
rect 324410 128616 324466 128625
rect 324410 128551 324466 128560
rect 324412 128308 324464 128314
rect 324412 128250 324464 128256
rect 324320 128240 324372 128246
rect 324320 128182 324372 128188
rect 324332 127809 324360 128182
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324424 127129 324452 128250
rect 324410 127120 324466 127129
rect 324410 127055 324466 127064
rect 324320 126948 324372 126954
rect 324320 126890 324372 126896
rect 324332 126313 324360 126890
rect 324318 126304 324374 126313
rect 324318 126239 324374 126248
rect 324516 125497 324544 132466
rect 324502 125488 324558 125497
rect 324502 125423 324558 125432
rect 325606 124808 325662 124817
rect 325712 124794 325740 210287
rect 325804 145489 325832 231066
rect 327080 219428 327132 219434
rect 327080 219370 327132 219376
rect 327092 219337 327120 219370
rect 327078 219328 327134 219337
rect 327078 219263 327134 219272
rect 327080 216028 327132 216034
rect 327080 215970 327132 215976
rect 325884 203584 325936 203590
rect 325884 203526 325936 203532
rect 325790 145480 325846 145489
rect 325790 145415 325846 145424
rect 325896 136377 325924 203526
rect 325974 177576 326030 177585
rect 325974 177511 326030 177520
rect 325988 170950 326016 177511
rect 325976 170944 326028 170950
rect 325976 170886 326028 170892
rect 325882 136368 325938 136377
rect 325882 136303 325938 136312
rect 325662 124766 325740 124794
rect 325606 124743 325662 124752
rect 324320 124160 324372 124166
rect 324320 124102 324372 124108
rect 324332 123185 324360 124102
rect 324318 123176 324374 123185
rect 324318 123111 324374 123120
rect 324320 122800 324372 122806
rect 324320 122742 324372 122748
rect 324332 122505 324360 122742
rect 324412 122732 324464 122738
rect 324412 122674 324464 122680
rect 324318 122496 324374 122505
rect 324318 122431 324374 122440
rect 324424 121689 324452 122674
rect 324410 121680 324466 121689
rect 324410 121615 324466 121624
rect 324412 121440 324464 121446
rect 324412 121382 324464 121388
rect 324320 121032 324372 121038
rect 324320 120974 324372 120980
rect 324332 120873 324360 120974
rect 324318 120864 324374 120873
rect 324318 120799 324374 120808
rect 324424 120193 324452 121382
rect 327092 121038 327120 215970
rect 327184 142089 327212 238002
rect 327276 209778 327304 434726
rect 328472 248414 328500 539582
rect 329840 499588 329892 499594
rect 329840 499530 329892 499536
rect 328472 248386 328592 248414
rect 328564 229022 328592 248386
rect 328552 229016 328604 229022
rect 328552 228958 328604 228964
rect 328564 227769 328592 228958
rect 328550 227760 328606 227769
rect 328550 227695 328606 227704
rect 329852 220833 329880 499530
rect 331496 354816 331548 354822
rect 331496 354758 331548 354764
rect 331312 239420 331364 239426
rect 331312 239362 331364 239368
rect 329932 227044 329984 227050
rect 329932 226986 329984 226992
rect 329838 220824 329894 220833
rect 329838 220759 329894 220768
rect 328460 214736 328512 214742
rect 328460 214678 328512 214684
rect 327264 209772 327316 209778
rect 327264 209714 327316 209720
rect 327276 209098 327304 209714
rect 327264 209092 327316 209098
rect 327264 209034 327316 209040
rect 327356 202156 327408 202162
rect 327356 202098 327408 202104
rect 327264 189780 327316 189786
rect 327264 189722 327316 189728
rect 327170 142080 327226 142089
rect 327170 142015 327226 142024
rect 327080 121032 327132 121038
rect 327080 120974 327132 120980
rect 324410 120184 324466 120193
rect 324410 120119 324466 120128
rect 324320 120080 324372 120086
rect 324320 120022 324372 120028
rect 324332 119377 324360 120022
rect 324318 119368 324374 119377
rect 324318 119303 324374 119312
rect 324412 118652 324464 118658
rect 324412 118594 324464 118600
rect 324320 118584 324372 118590
rect 324318 118552 324320 118561
rect 324372 118552 324374 118561
rect 324318 118487 324374 118496
rect 324424 117881 324452 118594
rect 324410 117872 324466 117881
rect 324410 117807 324466 117816
rect 323490 116512 323546 116521
rect 323490 116447 323546 116456
rect 323504 115977 323532 116447
rect 323490 115968 323546 115977
rect 323490 115903 323546 115912
rect 324412 115932 324464 115938
rect 324412 115874 324464 115880
rect 324320 115864 324372 115870
rect 324320 115806 324372 115812
rect 324332 115569 324360 115806
rect 324318 115560 324374 115569
rect 324318 115495 324374 115504
rect 324424 114753 324452 115874
rect 324410 114744 324466 114753
rect 324410 114679 324466 114688
rect 324320 114504 324372 114510
rect 324320 114446 324372 114452
rect 324332 114073 324360 114446
rect 324412 114436 324464 114442
rect 324412 114378 324464 114384
rect 324318 114064 324374 114073
rect 324318 113999 324374 114008
rect 324424 113257 324452 114378
rect 324410 113248 324466 113257
rect 324410 113183 324466 113192
rect 324320 113144 324372 113150
rect 324320 113086 324372 113092
rect 324332 112441 324360 113086
rect 324318 112432 324374 112441
rect 324318 112367 324374 112376
rect 324320 111784 324372 111790
rect 324318 111752 324320 111761
rect 324372 111752 324374 111761
rect 324318 111687 324374 111696
rect 324412 111716 324464 111722
rect 324412 111658 324464 111664
rect 324424 110945 324452 111658
rect 324410 110936 324466 110945
rect 324410 110871 324466 110880
rect 324320 110424 324372 110430
rect 324320 110366 324372 110372
rect 324332 110129 324360 110366
rect 324318 110120 324374 110129
rect 324318 110055 324374 110064
rect 323122 108624 323178 108633
rect 323122 108559 323178 108568
rect 323030 107128 323086 107137
rect 323030 107063 323086 107072
rect 322938 106312 322994 106321
rect 322938 106247 322994 106256
rect 321742 104272 321798 104281
rect 321742 104207 321798 104216
rect 321652 95124 321704 95130
rect 321652 95066 321704 95072
rect 321756 95062 321784 104207
rect 322938 100872 322994 100881
rect 322938 100807 322994 100816
rect 321834 98152 321890 98161
rect 321834 98087 321890 98096
rect 321744 95056 321796 95062
rect 321744 94998 321796 95004
rect 321560 93764 321612 93770
rect 321560 93706 321612 93712
rect 320180 90432 320232 90438
rect 320180 90374 320232 90380
rect 318064 78668 318116 78674
rect 318064 78610 318116 78616
rect 316132 76560 316184 76566
rect 316132 76502 316184 76508
rect 315304 75268 315356 75274
rect 315304 75210 315356 75216
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 309784 3460 309836 3466
rect 309784 3402 309836 3408
rect 310242 3360 310298 3369
rect 310242 3295 310298 3304
rect 310256 480 310284 3295
rect 311452 480 311480 16546
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 315316 4146 315344 75210
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 316144 3534 316172 76502
rect 317420 73704 317472 73710
rect 317420 73646 317472 73652
rect 317432 16574 317460 73646
rect 320192 16574 320220 90374
rect 321848 80034 321876 98087
rect 322952 81394 322980 100807
rect 323044 90982 323072 107063
rect 323136 95198 323164 108559
rect 324320 104848 324372 104854
rect 324320 104790 324372 104796
rect 324332 104009 324360 104790
rect 324318 104000 324374 104009
rect 324318 103935 324374 103944
rect 327276 103358 327304 189722
rect 327368 157214 327396 202098
rect 327356 157208 327408 157214
rect 327356 157150 327408 157156
rect 328472 104854 328500 214678
rect 328644 214600 328696 214606
rect 328644 214542 328696 214548
rect 328552 211880 328604 211886
rect 328552 211822 328604 211828
rect 328564 137902 328592 211822
rect 328656 151706 328684 214542
rect 329840 202292 329892 202298
rect 329840 202234 329892 202240
rect 328644 151700 328696 151706
rect 328644 151642 328696 151648
rect 328552 137896 328604 137902
rect 328552 137838 328604 137844
rect 329852 129742 329880 202234
rect 329840 129736 329892 129742
rect 329840 129678 329892 129684
rect 329944 128246 329972 226986
rect 330116 207732 330168 207738
rect 330116 207674 330168 207680
rect 330024 198008 330076 198014
rect 330024 197950 330076 197956
rect 330036 129674 330064 197950
rect 330128 154494 330156 207674
rect 331220 177472 331272 177478
rect 331220 177414 331272 177420
rect 331232 169726 331260 177414
rect 331220 169720 331272 169726
rect 331220 169662 331272 169668
rect 330116 154488 330168 154494
rect 330116 154430 330168 154436
rect 331324 133890 331352 239362
rect 331404 177540 331456 177546
rect 331404 177482 331456 177488
rect 331416 160070 331444 177482
rect 331404 160064 331456 160070
rect 331404 160006 331456 160012
rect 331312 133884 331364 133890
rect 331312 133826 331364 133832
rect 330024 129668 330076 129674
rect 330024 129610 330076 129616
rect 329932 128240 329984 128246
rect 329932 128182 329984 128188
rect 328460 104848 328512 104854
rect 328460 104790 328512 104796
rect 324320 103352 324372 103358
rect 324320 103294 324372 103300
rect 327264 103352 327316 103358
rect 327264 103294 327316 103300
rect 324332 103193 324360 103294
rect 324318 103184 324374 103193
rect 324318 103119 324374 103128
rect 324320 102128 324372 102134
rect 324320 102070 324372 102076
rect 324332 101697 324360 102070
rect 324318 101688 324374 101697
rect 324318 101623 324374 101632
rect 324502 100192 324558 100201
rect 324502 100127 324558 100136
rect 324410 99376 324466 99385
rect 324410 99311 324466 99320
rect 323124 95192 323176 95198
rect 323124 95134 323176 95140
rect 324424 93809 324452 99311
rect 324516 93838 324544 100127
rect 324594 97064 324650 97073
rect 324594 96999 324650 97008
rect 324504 93832 324556 93838
rect 324410 93800 324466 93809
rect 324504 93774 324556 93780
rect 324410 93735 324466 93744
rect 324608 92449 324636 96999
rect 324594 92440 324650 92449
rect 324594 92375 324650 92384
rect 323032 90976 323084 90982
rect 323032 90918 323084 90924
rect 328460 90364 328512 90370
rect 328460 90306 328512 90312
rect 324320 87712 324372 87718
rect 324320 87654 324372 87660
rect 323584 82136 323636 82142
rect 323584 82078 323636 82084
rect 322940 81388 322992 81394
rect 322940 81330 322992 81336
rect 321836 80028 321888 80034
rect 321836 79970 321888 79976
rect 317432 16546 318104 16574
rect 320192 16546 320496 16574
rect 316224 4140 316276 4146
rect 316224 4082 316276 4088
rect 316132 3528 316184 3534
rect 316132 3470 316184 3476
rect 315028 3188 315080 3194
rect 315028 3130 315080 3136
rect 315040 480 315068 3130
rect 316236 480 316264 4082
rect 317328 3528 317380 3534
rect 317328 3470 317380 3476
rect 317340 480 317368 3470
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319718 3632 319774 3641
rect 319718 3567 319774 3576
rect 319732 480 319760 3567
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 323596 3602 323624 82078
rect 323584 3596 323636 3602
rect 323584 3538 323636 3544
rect 322112 3460 322164 3466
rect 322112 3402 322164 3408
rect 322124 480 322152 3402
rect 324332 3346 324360 87654
rect 327080 82204 327132 82210
rect 327080 82146 327132 82152
rect 324412 25696 324464 25702
rect 324412 25638 324464 25644
rect 324424 3534 324452 25638
rect 327092 16574 327120 82146
rect 328472 16574 328500 90306
rect 331310 89040 331366 89049
rect 331310 88975 331366 88984
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 324412 3528 324464 3534
rect 324412 3470 324464 3476
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 323308 3324 323360 3330
rect 324332 3318 324452 3346
rect 323308 3266 323360 3272
rect 323320 480 323348 3266
rect 324424 480 324452 3318
rect 325620 480 325648 3470
rect 326804 3392 326856 3398
rect 326804 3334 326856 3340
rect 326816 480 326844 3334
rect 328012 480 328040 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330392 3256 330444 3262
rect 330392 3198 330444 3204
rect 330404 480 330432 3198
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331324 354 331352 88975
rect 331508 3262 331536 354758
rect 332612 230450 332640 565830
rect 332600 230444 332652 230450
rect 332600 230386 332652 230392
rect 332612 229094 332640 230386
rect 332612 229066 332732 229094
rect 332600 225616 332652 225622
rect 332600 225558 332652 225564
rect 332612 3534 332640 225558
rect 332704 186998 332732 229066
rect 333980 222896 334032 222902
rect 333980 222838 334032 222844
rect 332692 186992 332744 186998
rect 332692 186934 332744 186940
rect 332784 184408 332836 184414
rect 332784 184350 332836 184356
rect 332692 178764 332744 178770
rect 332692 178706 332744 178712
rect 332704 113150 332732 178706
rect 332796 158642 332824 184350
rect 332876 175976 332928 175982
rect 332876 175918 332928 175924
rect 332888 165510 332916 175918
rect 332876 165504 332928 165510
rect 332876 165446 332928 165452
rect 332784 158636 332836 158642
rect 332784 158578 332836 158584
rect 332692 113144 332744 113150
rect 332692 113086 332744 113092
rect 332690 21312 332746 21321
rect 332690 21247 332746 21256
rect 332600 3528 332652 3534
rect 332600 3470 332652 3476
rect 331496 3256 331548 3262
rect 331496 3198 331548 3204
rect 332704 480 332732 21247
rect 333992 16574 334020 222838
rect 335372 219434 335400 575486
rect 336004 320204 336056 320210
rect 336004 320146 336056 320152
rect 335452 232620 335504 232626
rect 335452 232562 335504 232568
rect 335360 219428 335412 219434
rect 335360 219370 335412 219376
rect 335360 210520 335412 210526
rect 335360 210462 335412 210468
rect 334256 195356 334308 195362
rect 334256 195298 334308 195304
rect 334072 181620 334124 181626
rect 334072 181562 334124 181568
rect 334084 111722 334112 181562
rect 334164 177336 334216 177342
rect 334164 177278 334216 177284
rect 334176 124166 334204 177278
rect 334268 164150 334296 195298
rect 335372 165578 335400 210462
rect 335360 165572 335412 165578
rect 335360 165514 335412 165520
rect 334256 164144 334308 164150
rect 334256 164086 334308 164092
rect 334164 124160 334216 124166
rect 334164 124102 334216 124108
rect 334072 111716 334124 111722
rect 334072 111658 334124 111664
rect 335464 16574 335492 232562
rect 335544 177404 335596 177410
rect 335544 177346 335596 177352
rect 335556 143546 335584 177346
rect 335544 143540 335596 143546
rect 335544 143482 335596 143488
rect 333992 16546 334664 16574
rect 335464 16546 335952 16574
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 333900 480 333928 3470
rect 331558 354 331670 480
rect 331324 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 335924 3482 335952 16546
rect 336016 4214 336044 320146
rect 336752 222057 336780 582354
rect 363616 549914 363644 696934
rect 363604 549908 363656 549914
rect 363604 549850 363656 549856
rect 349252 521688 349304 521694
rect 349252 521630 349304 521636
rect 347780 363724 347832 363730
rect 347780 363666 347832 363672
rect 337384 358828 337436 358834
rect 337384 358770 337436 358776
rect 336738 222048 336794 222057
rect 336738 221983 336794 221992
rect 336752 196761 336780 221983
rect 336738 196752 336794 196761
rect 336738 196687 336794 196696
rect 336922 184240 336978 184249
rect 336922 184175 336978 184184
rect 336832 182844 336884 182850
rect 336832 182786 336884 182792
rect 336740 181484 336792 181490
rect 336740 181426 336792 181432
rect 336752 115870 336780 181426
rect 336844 151774 336872 182786
rect 336936 157350 336964 184175
rect 336924 157344 336976 157350
rect 336924 157286 336976 157292
rect 336832 151768 336884 151774
rect 336832 151710 336884 151716
rect 336740 115864 336792 115870
rect 336740 115806 336792 115812
rect 336004 4208 336056 4214
rect 336004 4150 336056 4156
rect 335924 3454 336320 3482
rect 336292 480 336320 3454
rect 337396 2990 337424 358770
rect 342260 357536 342312 357542
rect 342260 357478 342312 357484
rect 339592 206304 339644 206310
rect 339592 206246 339644 206252
rect 339498 202192 339554 202201
rect 339498 202127 339554 202136
rect 338396 184272 338448 184278
rect 338396 184214 338448 184220
rect 338212 182980 338264 182986
rect 338212 182922 338264 182928
rect 338120 178696 338172 178702
rect 338120 178638 338172 178644
rect 338132 6186 338160 178638
rect 338224 139398 338252 182922
rect 338304 181688 338356 181694
rect 338304 181630 338356 181636
rect 338316 149054 338344 181630
rect 338408 168366 338436 184214
rect 338396 168360 338448 168366
rect 338396 168302 338448 168308
rect 338304 149048 338356 149054
rect 338304 148990 338356 148996
rect 338212 139392 338264 139398
rect 338212 139334 338264 139340
rect 339512 110430 339540 202127
rect 339604 118590 339632 206246
rect 340972 193860 341024 193866
rect 340972 193802 341024 193808
rect 340880 190052 340932 190058
rect 340880 189994 340932 190000
rect 339682 188320 339738 188329
rect 339682 188255 339738 188264
rect 339696 121446 339724 188255
rect 339776 184340 339828 184346
rect 339776 184282 339828 184288
rect 339788 164218 339816 184282
rect 339776 164212 339828 164218
rect 339776 164154 339828 164160
rect 339684 121440 339736 121446
rect 339684 121382 339736 121388
rect 339592 118584 339644 118590
rect 339592 118526 339644 118532
rect 339500 110424 339552 110430
rect 339500 110366 339552 110372
rect 338120 6180 338172 6186
rect 338120 6122 338172 6128
rect 337476 3596 337528 3602
rect 337476 3538 337528 3544
rect 337384 2984 337436 2990
rect 337384 2926 337436 2932
rect 337488 480 337516 3538
rect 340892 3534 340920 189994
rect 340984 120086 341012 193802
rect 341064 189848 341116 189854
rect 341064 189790 341116 189796
rect 341076 161430 341104 189790
rect 341156 180124 341208 180130
rect 341156 180066 341208 180072
rect 341064 161424 341116 161430
rect 341064 161366 341116 161372
rect 341168 153202 341196 180066
rect 341156 153196 341208 153202
rect 341156 153138 341208 153144
rect 340972 120080 341024 120086
rect 340972 120022 341024 120028
rect 340972 4208 341024 4214
rect 340972 4150 341024 4156
rect 340880 3528 340932 3534
rect 340880 3470 340932 3476
rect 338672 2984 338724 2990
rect 338672 2926 338724 2932
rect 338684 480 338712 2926
rect 339866 2000 339922 2009
rect 339866 1935 339922 1944
rect 339880 480 339908 1935
rect 340984 480 341012 4150
rect 342166 3496 342222 3505
rect 342166 3431 342222 3440
rect 342180 480 342208 3431
rect 342272 3330 342300 357478
rect 345664 356176 345716 356182
rect 345664 356118 345716 356124
rect 343640 221468 343692 221474
rect 343640 221410 343692 221416
rect 342352 203652 342404 203658
rect 342352 203594 342404 203600
rect 342364 16574 342392 203594
rect 342442 200696 342498 200705
rect 342442 200631 342498 200640
rect 342456 135182 342484 200631
rect 342536 191208 342588 191214
rect 342536 191150 342588 191156
rect 342444 135176 342496 135182
rect 342444 135118 342496 135124
rect 342548 126954 342576 191150
rect 342628 179308 342680 179314
rect 342628 179250 342680 179256
rect 342640 179217 342668 179250
rect 342626 179208 342682 179217
rect 342626 179143 342682 179152
rect 342536 126948 342588 126954
rect 342536 126890 342588 126896
rect 343652 114442 343680 221410
rect 345020 206508 345072 206514
rect 345020 206450 345072 206456
rect 343732 204944 343784 204950
rect 343732 204886 343784 204892
rect 343744 122738 343772 204886
rect 343914 180024 343970 180033
rect 343914 179959 343970 179968
rect 343824 175296 343876 175302
rect 343824 175238 343876 175244
rect 343836 131102 343864 175238
rect 343928 158710 343956 179959
rect 343916 158704 343968 158710
rect 343916 158646 343968 158652
rect 343824 131096 343876 131102
rect 343824 131038 343876 131044
rect 343732 122732 343784 122738
rect 343732 122674 343784 122680
rect 343640 114436 343692 114442
rect 343640 114378 343692 114384
rect 345032 111790 345060 206450
rect 345204 182912 345256 182918
rect 345204 182854 345256 182860
rect 345112 181552 345164 181558
rect 345112 181494 345164 181500
rect 345124 137970 345152 181494
rect 345216 144906 345244 182854
rect 345204 144900 345256 144906
rect 345204 144842 345256 144848
rect 345112 137964 345164 137970
rect 345112 137906 345164 137912
rect 345020 111784 345072 111790
rect 345020 111726 345072 111732
rect 345676 33114 345704 356118
rect 347044 327752 347096 327758
rect 347044 327694 347096 327700
rect 347056 259418 347084 327694
rect 347044 259412 347096 259418
rect 347044 259354 347096 259360
rect 347044 242956 347096 242962
rect 347044 242898 347096 242904
rect 347056 233238 347084 242898
rect 347044 233232 347096 233238
rect 347044 233174 347096 233180
rect 346584 231872 346636 231878
rect 346584 231814 346636 231820
rect 346492 205080 346544 205086
rect 346492 205022 346544 205028
rect 346400 192772 346452 192778
rect 346400 192714 346452 192720
rect 346308 179376 346360 179382
rect 346306 179344 346308 179353
rect 346360 179344 346362 179353
rect 346306 179279 346362 179288
rect 345664 33108 345716 33114
rect 345664 33050 345716 33056
rect 343640 32496 343692 32502
rect 343640 32438 343692 32444
rect 343652 16574 343680 32438
rect 345662 18728 345718 18737
rect 345662 18663 345718 18672
rect 345020 17400 345072 17406
rect 345020 17342 345072 17348
rect 345032 16574 345060 17342
rect 342364 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 342260 3324 342312 3330
rect 342260 3266 342312 3272
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 345676 3194 345704 18663
rect 346412 16574 346440 192714
rect 346504 114510 346532 205022
rect 346596 154562 346624 231814
rect 346676 216708 346728 216714
rect 346676 216650 346728 216656
rect 346584 154556 346636 154562
rect 346584 154498 346636 154504
rect 346688 150414 346716 216650
rect 346676 150408 346728 150414
rect 346676 150350 346728 150356
rect 347792 147626 347820 363666
rect 349264 234598 349292 521630
rect 364352 472666 364380 702406
rect 397472 699718 397500 703520
rect 413664 702642 413692 703520
rect 413652 702636 413704 702642
rect 413652 702578 413704 702584
rect 395344 699712 395396 699718
rect 395344 699654 395396 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 364340 472660 364392 472666
rect 364340 472602 364392 472608
rect 353300 392012 353352 392018
rect 353300 391954 353352 391960
rect 350540 318844 350592 318850
rect 350540 318786 350592 318792
rect 349344 269136 349396 269142
rect 349344 269078 349396 269084
rect 349252 234592 349304 234598
rect 349252 234534 349304 234540
rect 347872 199436 347924 199442
rect 347872 199378 347924 199384
rect 347780 147620 347832 147626
rect 347780 147562 347832 147568
rect 347884 118658 347912 199378
rect 347964 184204 348016 184210
rect 347964 184146 348016 184152
rect 347976 128314 348004 184146
rect 347964 128308 348016 128314
rect 347964 128250 348016 128256
rect 347872 118652 347924 118658
rect 347872 118594 347924 118600
rect 346492 114504 346544 114510
rect 346492 114446 346544 114452
rect 349264 102134 349292 234534
rect 349252 102128 349304 102134
rect 349252 102070 349304 102076
rect 347778 50280 347834 50289
rect 347778 50215 347834 50224
rect 347792 16574 347820 50215
rect 349356 16574 349384 269078
rect 350552 16574 350580 318786
rect 350632 206372 350684 206378
rect 350632 206314 350684 206320
rect 350644 135250 350672 206314
rect 351920 200796 351972 200802
rect 351920 200738 351972 200744
rect 350632 135244 350684 135250
rect 350632 135186 350684 135192
rect 351932 122806 351960 200738
rect 353312 162858 353340 391954
rect 395356 375329 395384 699654
rect 429856 698970 429884 703520
rect 462332 702574 462360 703520
rect 462320 702568 462372 702574
rect 462320 702510 462372 702516
rect 478524 702434 478552 703520
rect 494808 702778 494836 703520
rect 494796 702772 494848 702778
rect 494796 702714 494848 702720
rect 527192 702710 527220 703520
rect 527180 702704 527232 702710
rect 527180 702646 527232 702652
rect 543476 702506 543504 703520
rect 543464 702500 543516 702506
rect 543464 702442 543516 702448
rect 477512 702406 478552 702434
rect 429844 698964 429896 698970
rect 429844 698906 429896 698912
rect 445024 563100 445076 563106
rect 445024 563042 445076 563048
rect 445036 404326 445064 563042
rect 445024 404320 445076 404326
rect 445024 404262 445076 404268
rect 477512 400178 477540 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580262 617536 580318 617545
rect 580262 617471 580318 617480
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 589966 580212 590951
rect 580172 589960 580224 589966
rect 580172 589902 580224 589908
rect 579804 578196 579856 578202
rect 579804 578138 579856 578144
rect 579816 577697 579844 578138
rect 579802 577688 579858 577697
rect 579802 577623 579858 577632
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 500224 556232 500276 556238
rect 500224 556174 500276 556180
rect 500236 419490 500264 556174
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580276 482322 580304 617471
rect 580354 524512 580410 524521
rect 580354 524447 580410 524456
rect 580264 482316 580316 482322
rect 580264 482258 580316 482264
rect 580078 471472 580134 471481
rect 580078 471407 580134 471416
rect 580092 470626 580120 471407
rect 580080 470620 580132 470626
rect 580080 470562 580132 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 500224 419484 500276 419490
rect 500224 419426 500276 419432
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580368 407794 580396 524447
rect 582378 431624 582434 431633
rect 582378 431559 582434 431568
rect 580356 407788 580408 407794
rect 580356 407730 580408 407736
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 477500 400172 477552 400178
rect 477500 400114 477552 400120
rect 582392 396778 582420 431559
rect 582380 396772 582432 396778
rect 582380 396714 582432 396720
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 395342 375320 395398 375329
rect 395342 375255 395398 375264
rect 356060 372632 356112 372638
rect 356060 372574 356112 372580
rect 355324 309800 355376 309806
rect 355324 309742 355376 309748
rect 353944 235272 353996 235278
rect 353944 235214 353996 235220
rect 353300 162852 353352 162858
rect 353300 162794 353352 162800
rect 351920 122800 351972 122806
rect 351920 122742 351972 122748
rect 353956 46918 353984 235214
rect 355336 219434 355364 309742
rect 355324 219428 355376 219434
rect 355324 219370 355376 219376
rect 354680 209092 354732 209098
rect 354680 209034 354732 209040
rect 354692 115938 354720 209034
rect 354772 196852 354824 196858
rect 354772 196794 354824 196800
rect 354784 132462 354812 196794
rect 356072 155922 356100 372574
rect 580906 365120 580962 365129
rect 580906 365055 580962 365064
rect 580920 363662 580948 365055
rect 582380 364404 582432 364410
rect 582380 364346 582432 364352
rect 580908 363656 580960 363662
rect 580908 363598 580960 363604
rect 580264 360256 580316 360262
rect 580264 360198 580316 360204
rect 449164 357468 449216 357474
rect 449164 357410 449216 357416
rect 356704 313336 356756 313342
rect 356704 313278 356756 313284
rect 356060 155916 356112 155922
rect 356060 155858 356112 155864
rect 354772 132456 354824 132462
rect 354772 132398 354824 132404
rect 354680 115932 354732 115938
rect 354680 115874 354732 115880
rect 356716 73166 356744 313278
rect 359464 281580 359516 281586
rect 359464 281522 359516 281528
rect 356704 73160 356756 73166
rect 356704 73102 356756 73108
rect 359476 60722 359504 281522
rect 449176 126954 449204 357410
rect 580276 351937 580304 360198
rect 580262 351928 580318 351937
rect 580262 351863 580318 351872
rect 468484 345704 468536 345710
rect 468484 345646 468536 345652
rect 467104 316736 467156 316742
rect 467104 316678 467156 316684
rect 449164 126948 449216 126954
rect 449164 126890 449216 126896
rect 467116 113150 467144 316678
rect 468496 139398 468524 345646
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 512644 245676 512696 245682
rect 512644 245618 512696 245624
rect 468484 139392 468536 139398
rect 468484 139334 468536 139340
rect 467104 113144 467156 113150
rect 467104 113086 467156 113092
rect 512656 100706 512684 245618
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 240106 580212 245511
rect 580262 240816 580318 240825
rect 580262 240751 580318 240760
rect 580172 240100 580224 240106
rect 580172 240042 580224 240048
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 574744 229764 574796 229770
rect 574744 229706 574796 229712
rect 574756 206990 574784 229706
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 574744 206984 574796 206990
rect 574744 206926 574796 206932
rect 579896 206984 579948 206990
rect 579896 206926 579948 206932
rect 579908 205737 579936 206926
rect 579894 205728 579950 205737
rect 579894 205663 579950 205672
rect 580276 179217 580304 240751
rect 580354 226944 580410 226953
rect 580354 226879 580410 226888
rect 580368 192545 580396 226879
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 580262 179208 580318 179217
rect 580262 179143 580318 179152
rect 582392 152697 582420 364346
rect 582562 354512 582618 354521
rect 582562 354447 582618 354456
rect 582470 272232 582526 272241
rect 582470 272167 582526 272176
rect 582484 238649 582512 272167
rect 582470 238640 582526 238649
rect 582470 238575 582526 238584
rect 582472 195288 582524 195294
rect 582472 195230 582524 195236
rect 582378 152688 582434 152697
rect 582378 152623 582434 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 512644 100700 512696 100706
rect 512644 100642 512696 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 359464 60716 359516 60722
rect 359464 60658 359516 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 353944 46912 353996 46918
rect 353944 46854 353996 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579618 39264 579674 39273
rect 579618 39199 579674 39208
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 349356 16546 350488 16574
rect 350552 16546 351224 16574
rect 345664 3188 345716 3194
rect 345664 3130 345716 3136
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349252 3188 349304 3194
rect 349252 3130 349304 3136
rect 349264 480 349292 3130
rect 350460 480 350488 16546
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579632 354 579660 39199
rect 579894 33144 579950 33153
rect 579894 33079 579896 33088
rect 579948 33079 579950 33088
rect 579896 33050 579948 33056
rect 579896 20664 579948 20670
rect 579896 20606 579948 20612
rect 579908 19825 579936 20606
rect 579894 19816 579950 19825
rect 579894 19751 579950 19760
rect 582484 6633 582512 195230
rect 582576 165889 582604 354447
rect 582562 165880 582618 165889
rect 582562 165815 582618 165824
rect 582470 6624 582526 6633
rect 582470 6559 582526 6568
rect 579774 354 579886 480
rect 579632 326 579886 354
rect 579774 -960 579886 326
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 606076 3570 606112
rect 3514 606056 3516 606076
rect 3516 606056 3568 606076
rect 3568 606056 3570 606076
rect 2870 579944 2926 580000
rect 3422 566888 3478 566944
rect 3146 553832 3202 553888
rect 3698 527856 3754 527912
rect 3422 514800 3478 514856
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3422 462576 3478 462632
rect 3330 449520 3386 449576
rect 3422 423544 3478 423600
rect 3422 410488 3478 410544
rect 3974 397432 4030 397488
rect 3422 371320 3478 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 1306 177248 1362 177304
rect 2870 293120 2926 293176
rect 3422 267144 3478 267200
rect 3422 254088 3478 254144
rect 2962 241032 3018 241088
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 2778 162832 2834 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3514 84632 3570 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 2778 37848 2834 37904
rect 2686 16496 2742 16552
rect 1398 15272 1454 15328
rect 2686 15272 2742 15328
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 16578 62736 16634 62792
rect 13818 59880 13874 59936
rect 3422 6432 3478 6488
rect 31666 558184 31722 558240
rect 27618 18536 27674 18592
rect 30102 12960 30158 13016
rect 37186 301416 37242 301472
rect 41326 586336 41382 586392
rect 39854 357992 39910 358048
rect 39854 284280 39910 284336
rect 44086 403688 44142 403744
rect 35898 48864 35954 48920
rect 49514 341400 49570 341456
rect 50986 585248 51042 585304
rect 52366 401648 52422 401704
rect 53562 405592 53618 405648
rect 53746 464888 53802 464944
rect 54942 403552 54998 403608
rect 53838 284300 53894 284336
rect 53838 284280 53840 284300
rect 53840 284280 53892 284300
rect 53892 284280 53894 284300
rect 52182 200776 52238 200832
rect 54942 271768 54998 271824
rect 54850 225528 54906 225584
rect 58622 586608 58678 586664
rect 57794 583752 57850 583808
rect 56230 238720 56286 238776
rect 58622 469784 58678 469840
rect 58714 434560 58770 434616
rect 59174 314744 59230 314800
rect 57702 202272 57758 202328
rect 52550 177248 52606 177304
rect 52458 58520 52514 58576
rect 52550 26832 52606 26888
rect 61382 585112 61438 585168
rect 60738 568928 60794 568984
rect 60738 565528 60794 565584
rect 60738 562128 60794 562184
rect 60738 555328 60794 555384
rect 60738 552608 60794 552664
rect 60738 549208 60794 549264
rect 60738 542428 60794 542464
rect 60738 542408 60740 542428
rect 60740 542408 60792 542428
rect 60792 542408 60794 542428
rect 60738 539008 60794 539064
rect 60738 535608 60794 535664
rect 60738 528808 60794 528864
rect 60370 518608 60426 518664
rect 60738 515208 60794 515264
rect 60554 505008 60610 505064
rect 60738 502288 60794 502344
rect 60738 495508 60794 495544
rect 60738 495488 60740 495508
rect 60740 495488 60792 495508
rect 60792 495488 60794 495508
rect 60738 492088 60794 492144
rect 61658 522008 61714 522064
rect 62026 545808 62082 545864
rect 61934 510448 61990 510504
rect 61934 508408 61990 508464
rect 60738 488688 60794 488744
rect 61842 485832 61898 485888
rect 61198 485288 61254 485344
rect 61566 481888 61622 481944
rect 60738 478488 60794 478544
rect 61382 475088 61438 475144
rect 60922 471688 60978 471744
rect 60738 468288 60794 468344
rect 60738 464888 60794 464944
rect 60738 461488 60794 461544
rect 60738 458088 60794 458144
rect 61842 473184 61898 473240
rect 61750 454688 61806 454744
rect 60738 445168 60794 445224
rect 60738 441768 60794 441824
rect 60922 438368 60978 438424
rect 61566 434968 61622 435024
rect 60738 428168 60794 428224
rect 60738 424768 60794 424824
rect 60738 414568 60794 414624
rect 60738 407788 60794 407824
rect 60738 407768 60740 407788
rect 60740 407768 60792 407788
rect 60792 407768 60794 407788
rect 61842 451968 61898 452024
rect 61842 359352 61898 359408
rect 61750 239400 61806 239456
rect 62302 417968 62358 418024
rect 63038 498888 63094 498944
rect 63314 525408 63370 525464
rect 63314 449928 63370 449984
rect 83370 586608 83426 586664
rect 99378 586336 99434 586392
rect 169666 585384 169722 585440
rect 178682 585248 178738 585304
rect 201406 586336 201462 586392
rect 232778 586608 232834 586664
rect 64418 584568 64474 584624
rect 92754 584568 92810 584624
rect 188066 584568 188122 584624
rect 223486 584568 223542 584624
rect 243266 585112 243322 585168
rect 243634 585112 243690 585168
rect 243542 580896 243598 580952
rect 63498 471688 63554 471744
rect 63406 438368 63462 438424
rect 63222 429256 63278 429312
rect 63682 410624 63738 410680
rect 63130 253952 63186 254008
rect 63406 252456 63462 252512
rect 242806 405456 242862 405512
rect 66166 404504 66222 404560
rect 65522 404368 65578 404424
rect 64694 294480 64750 294536
rect 67638 399472 67694 399528
rect 67546 296792 67602 296848
rect 67730 291080 67786 291136
rect 67638 290400 67694 290456
rect 67730 289720 67786 289776
rect 67638 289040 67694 289096
rect 67638 287680 67694 287736
rect 67822 287000 67878 287056
rect 67730 286320 67786 286376
rect 67638 284316 67640 284336
rect 67640 284316 67692 284336
rect 67692 284316 67694 284336
rect 67638 284280 67694 284316
rect 67730 283600 67786 283656
rect 67638 282920 67694 282976
rect 68742 292848 68798 292904
rect 68742 284960 68798 285016
rect 68650 281560 68706 281616
rect 67638 280880 67694 280936
rect 67638 280220 67694 280256
rect 67638 280200 67640 280220
rect 67640 280200 67692 280220
rect 67692 280200 67694 280220
rect 67638 279520 67694 279576
rect 67730 278840 67786 278896
rect 67638 278160 67694 278216
rect 67638 277480 67694 277536
rect 69110 285640 69166 285696
rect 67730 276800 67786 276856
rect 67638 276140 67694 276176
rect 67638 276120 67640 276140
rect 67640 276120 67692 276140
rect 67692 276120 67694 276140
rect 68190 275476 68192 275496
rect 68192 275476 68244 275496
rect 68244 275476 68246 275496
rect 68190 275440 68246 275476
rect 67638 274760 67694 274816
rect 68006 274080 68062 274136
rect 67822 273400 67878 273456
rect 67638 272720 67694 272776
rect 67822 272040 67878 272096
rect 67730 271360 67786 271416
rect 67638 270680 67694 270736
rect 67730 270000 67786 270056
rect 67638 269320 67694 269376
rect 67730 268640 67786 268696
rect 67638 267960 67694 268016
rect 68926 275440 68982 275496
rect 68650 267280 68706 267336
rect 67546 266600 67602 266656
rect 68098 265920 68154 265976
rect 67638 265240 67694 265296
rect 67638 264560 67694 264616
rect 68834 263880 68890 263936
rect 67730 263200 67786 263256
rect 67638 262520 67694 262576
rect 67638 261840 67694 261896
rect 67730 261160 67786 261216
rect 67638 260480 67694 260536
rect 67730 259800 67786 259856
rect 67730 259120 67786 259176
rect 67638 258440 67694 258496
rect 67638 257760 67694 257816
rect 67638 256400 67694 256456
rect 67914 255720 67970 255776
rect 68742 255720 68798 255776
rect 67730 255040 67786 255096
rect 67638 254360 67694 254416
rect 67638 253680 67694 253736
rect 67638 251640 67694 251696
rect 67638 250960 67694 251016
rect 67546 250280 67602 250336
rect 66902 238448 66958 238504
rect 67638 249600 67694 249656
rect 67638 248920 67694 248976
rect 67730 248240 67786 248296
rect 67638 247560 67694 247616
rect 67638 246880 67694 246936
rect 68190 246200 68246 246256
rect 68190 244840 68246 244896
rect 67638 243480 67694 243536
rect 67638 242800 67694 242856
rect 67730 242120 67786 242176
rect 67638 241460 67694 241496
rect 67638 241440 67640 241460
rect 67640 241440 67692 241460
rect 67692 241440 67694 241460
rect 67638 240760 67694 240816
rect 69110 274080 69166 274136
rect 70490 292304 70546 292360
rect 71778 295316 71834 295352
rect 71778 295296 71780 295316
rect 71780 295296 71832 295316
rect 71832 295296 71834 295316
rect 73158 404912 73214 404968
rect 76010 398112 76066 398168
rect 73710 301144 73766 301200
rect 73894 295160 73950 295216
rect 75826 294480 75882 294536
rect 76010 294480 76066 294536
rect 78402 294208 78458 294264
rect 90362 397976 90418 398032
rect 89718 304952 89774 305008
rect 90362 304952 90418 305008
rect 88982 303612 89038 303648
rect 88982 303592 88984 303612
rect 88984 303592 89036 303612
rect 89036 303592 89038 303612
rect 95882 380160 95938 380216
rect 103518 403552 103574 403608
rect 103426 296928 103482 296984
rect 103518 295432 103574 295488
rect 108946 389816 109002 389872
rect 105542 386960 105598 387016
rect 104346 296928 104402 296984
rect 104162 295432 104218 295488
rect 105542 292712 105598 292768
rect 106094 292712 106150 292768
rect 107658 300736 107714 300792
rect 108946 300736 109002 300792
rect 108946 299512 109002 299568
rect 110326 349696 110382 349752
rect 109130 301008 109186 301064
rect 110326 301008 110382 301064
rect 113178 354728 113234 354784
rect 112442 298832 112498 298888
rect 111890 294072 111946 294128
rect 113822 292576 113878 292632
rect 118606 400832 118662 400888
rect 117686 295568 117742 295624
rect 118974 298832 119030 298888
rect 118606 295568 118662 295624
rect 117962 292032 118018 292088
rect 119066 291896 119122 291952
rect 69202 265920 69258 265976
rect 120078 286320 120134 286376
rect 120170 280880 120226 280936
rect 69662 243616 69718 243672
rect 120170 250960 120226 251016
rect 120630 250960 120686 251016
rect 119894 240896 119950 240952
rect 72606 238584 72662 238640
rect 72606 237088 72662 237144
rect 74538 238720 74594 238776
rect 86130 238584 86186 238640
rect 85486 222808 85542 222864
rect 80702 185544 80758 185600
rect 109038 238720 109094 238776
rect 109958 238720 110014 238776
rect 111154 239264 111210 239320
rect 68926 181328 68982 181384
rect 100666 177520 100722 177576
rect 102046 177520 102102 177576
rect 104806 177520 104862 177576
rect 106186 177520 106242 177576
rect 107014 176740 107016 176760
rect 107016 176740 107068 176760
rect 107068 176740 107070 176760
rect 107014 176704 107070 176740
rect 108118 176704 108174 176760
rect 109958 176704 110014 176760
rect 114466 236952 114522 237008
rect 117686 238468 117742 238504
rect 117686 238448 117688 238468
rect 117688 238448 117740 238468
rect 117740 238448 117742 238468
rect 120078 241440 120134 241496
rect 117962 195200 118018 195256
rect 114006 182144 114062 182200
rect 114006 177520 114062 177576
rect 121458 291760 121514 291816
rect 121458 290400 121514 290456
rect 121458 289040 121514 289096
rect 121458 287680 121514 287736
rect 121642 291080 121698 291136
rect 121642 288360 121698 288416
rect 121458 284960 121514 285016
rect 121550 284280 121606 284336
rect 121458 282940 121514 282976
rect 121458 282920 121460 282940
rect 121460 282920 121512 282940
rect 121512 282920 121514 282940
rect 121550 282240 121606 282296
rect 121458 281580 121514 281616
rect 121458 281560 121460 281580
rect 121460 281560 121512 281580
rect 121512 281560 121514 281580
rect 121458 280220 121514 280256
rect 121458 280200 121460 280220
rect 121460 280200 121512 280220
rect 121512 280200 121514 280220
rect 121458 278840 121514 278896
rect 122102 280880 122158 280936
rect 121642 278704 121698 278760
rect 121550 277480 121606 277536
rect 121458 276800 121514 276856
rect 121458 275440 121514 275496
rect 121550 274760 121606 274816
rect 121458 274080 121514 274136
rect 121458 273400 121514 273456
rect 121458 272720 121514 272776
rect 121458 271360 121514 271416
rect 121458 270000 121514 270056
rect 121550 269320 121606 269376
rect 121458 268640 121514 268696
rect 121458 267960 121514 268016
rect 121458 267280 121514 267336
rect 121550 266600 121606 266656
rect 121458 264560 121514 264616
rect 121550 263880 121606 263936
rect 121458 263200 121514 263256
rect 121458 262520 121514 262576
rect 120998 261840 121054 261896
rect 121458 261160 121514 261216
rect 121458 260480 121514 260536
rect 122746 279520 122802 279576
rect 122286 278704 122342 278760
rect 122194 265920 122250 265976
rect 121458 259800 121514 259856
rect 122102 259120 122158 259176
rect 121458 258440 121514 258496
rect 121550 257760 121606 257816
rect 121458 257080 121514 257136
rect 121550 256400 121606 256456
rect 121458 255720 121514 255776
rect 121458 254360 121514 254416
rect 121550 253680 121606 253736
rect 121458 253000 121514 253056
rect 121458 252320 121514 252376
rect 121550 250280 121606 250336
rect 121458 249600 121514 249656
rect 121550 248240 121606 248296
rect 121458 247560 121514 247616
rect 121550 246880 121606 246936
rect 121458 246200 121514 246256
rect 121458 245520 121514 245576
rect 121550 244840 121606 244896
rect 121458 244196 121460 244216
rect 121460 244196 121512 244216
rect 121512 244196 121514 244216
rect 121458 244160 121514 244196
rect 121458 242820 121514 242856
rect 121458 242800 121460 242820
rect 121460 242800 121512 242820
rect 121512 242800 121514 242820
rect 121550 242120 121606 242176
rect 121458 240760 121514 240816
rect 121550 240080 121606 240136
rect 122378 272040 122434 272096
rect 122194 251640 122250 251696
rect 122102 228928 122158 228984
rect 122378 255040 122434 255096
rect 122930 248920 122986 248976
rect 124402 286592 124458 286648
rect 126886 341400 126942 341456
rect 128358 240896 128414 240952
rect 131026 362208 131082 362264
rect 129186 204856 129242 204912
rect 118422 177520 118478 177576
rect 122010 177520 122066 177576
rect 132590 356088 132646 356144
rect 130382 181600 130438 181656
rect 125506 177520 125562 177576
rect 114282 176976 114338 177032
rect 120998 176976 121054 177032
rect 123022 176976 123078 177032
rect 139490 327664 139546 327720
rect 141514 294072 141570 294128
rect 142802 291896 142858 291952
rect 143630 301416 143686 301472
rect 145746 272584 145802 272640
rect 147586 400968 147642 401024
rect 149058 298696 149114 298752
rect 147586 266192 147642 266248
rect 147586 265512 147642 265568
rect 147126 241168 147182 241224
rect 142802 188400 142858 188456
rect 151818 376624 151874 376680
rect 152554 376624 152610 376680
rect 152554 375400 152610 375456
rect 149886 193976 149942 194032
rect 151082 186904 151138 186960
rect 151174 182824 151230 182880
rect 132406 177520 132462 177576
rect 133602 177520 133658 177576
rect 112442 176704 112498 176760
rect 125782 176704 125838 176760
rect 127070 176704 127126 176760
rect 128174 176704 128230 176760
rect 130750 176704 130806 176760
rect 134430 176704 134486 176760
rect 135718 176724 135774 176760
rect 135718 176704 135720 176724
rect 135720 176704 135772 176724
rect 135772 176704 135774 176724
rect 148230 176704 148286 176760
rect 98366 175344 98422 175400
rect 100758 175344 100814 175400
rect 116950 175344 117006 175400
rect 152646 190984 152702 191040
rect 159362 403552 159418 403608
rect 157982 296792 158038 296848
rect 158626 238584 158682 238640
rect 158626 237360 158682 237416
rect 161754 357992 161810 358048
rect 161478 357448 161534 357504
rect 161754 357448 161810 357504
rect 160742 237360 160798 237416
rect 162766 314744 162822 314800
rect 161478 224168 161534 224224
rect 162214 298696 162270 298752
rect 163502 237224 163558 237280
rect 164238 353368 164294 353424
rect 165434 354592 165490 354648
rect 165434 353368 165490 353424
rect 162306 192480 162362 192536
rect 162122 178608 162178 178664
rect 159914 176704 159970 176760
rect 165526 241440 165582 241496
rect 165526 240760 165582 240816
rect 164882 181464 164938 181520
rect 162398 176568 162454 176624
rect 152554 175888 152610 175944
rect 129462 175344 129518 175400
rect 115754 174936 115810 174992
rect 119434 174936 119490 174992
rect 67546 129240 67602 129296
rect 66166 128016 66222 128072
rect 64786 127064 64842 127120
rect 66166 127064 66222 127120
rect 64694 102176 64750 102232
rect 66166 126248 66222 126304
rect 66166 125160 66222 125216
rect 66074 122576 66130 122632
rect 67454 123528 67510 123584
rect 67362 120808 67418 120864
rect 67638 100680 67694 100736
rect 67546 94832 67602 94888
rect 67454 89664 67510 89720
rect 166998 290400 167054 290456
rect 167826 294208 167882 294264
rect 167826 238720 167882 238776
rect 166906 177248 166962 177304
rect 166538 176568 166594 176624
rect 169114 292848 169170 292904
rect 169298 292712 169354 292768
rect 170770 231784 170826 231840
rect 167918 171536 167974 171592
rect 109038 94696 109094 94752
rect 113730 94696 113786 94752
rect 131946 94696 132002 94752
rect 151726 94696 151782 94752
rect 151910 94696 151966 94752
rect 121734 93608 121790 93664
rect 102046 93472 102102 93528
rect 107750 93472 107806 93528
rect 124494 93472 124550 93528
rect 110142 93200 110198 93256
rect 119342 93200 119398 93256
rect 74814 92384 74870 92440
rect 85946 92384 86002 92440
rect 94226 92384 94282 92440
rect 101862 92384 101918 92440
rect 85026 91160 85082 91216
rect 89074 91704 89130 91760
rect 86774 91160 86830 91216
rect 87418 91160 87474 91216
rect 99286 91432 99342 91488
rect 97906 91296 97962 91352
rect 99102 91296 99158 91352
rect 91006 91160 91062 91216
rect 92386 91160 92442 91216
rect 93766 91160 93822 91216
rect 95054 91160 95110 91216
rect 96526 91160 96582 91216
rect 97814 91160 97870 91216
rect 56598 8880 56654 8936
rect 99194 91160 99250 91216
rect 99194 78512 99250 78568
rect 104530 91568 104586 91624
rect 106922 91568 106978 91624
rect 99930 91160 99986 91216
rect 100666 91160 100722 91216
rect 102046 91160 102102 91216
rect 102966 91160 103022 91216
rect 103426 91160 103482 91216
rect 104622 91160 104678 91216
rect 106186 91160 106242 91216
rect 106646 91160 106702 91216
rect 104622 86808 104678 86864
rect 115202 92384 115258 92440
rect 115478 92384 115534 92440
rect 120354 92404 120410 92440
rect 120354 92384 120356 92404
rect 120356 92384 120408 92404
rect 120408 92384 120410 92404
rect 112350 91704 112406 91760
rect 110326 91160 110382 91216
rect 110694 91160 110750 91216
rect 111706 91160 111762 91216
rect 110694 88168 110750 88224
rect 110326 84088 110382 84144
rect 114466 91160 114522 91216
rect 124126 92384 124182 92440
rect 125966 92384 126022 92440
rect 133142 92384 133198 92440
rect 151726 92384 151782 92440
rect 123942 91704 123998 91760
rect 122838 91432 122894 91488
rect 118238 91296 118294 91352
rect 115754 91160 115810 91216
rect 116766 91160 116822 91216
rect 117134 91160 117190 91216
rect 118606 91160 118662 91216
rect 119986 91160 120042 91216
rect 121090 91160 121146 91216
rect 122378 91160 122434 91216
rect 151726 91704 151782 91760
rect 126610 91568 126666 91624
rect 125506 91160 125562 91216
rect 126886 91160 126942 91216
rect 88338 69536 88394 69592
rect 129646 91160 129702 91216
rect 131026 91160 131082 91216
rect 135074 91160 135130 91216
rect 135902 91160 135958 91216
rect 166262 88168 166318 88224
rect 167918 111732 167920 111752
rect 167920 111732 167972 111752
rect 167972 111732 167974 111752
rect 167918 111696 167974 111732
rect 168102 110064 168158 110120
rect 167918 108704 167974 108760
rect 171874 295296 171930 295352
rect 172426 295296 172482 295352
rect 173714 293936 173770 293992
rect 172334 255176 172390 255232
rect 176566 403688 176622 403744
rect 172058 93880 172114 93936
rect 173346 92112 173402 92168
rect 125874 3304 125930 3360
rect 176658 354356 176660 354376
rect 176660 354356 176712 354376
rect 176712 354356 176714 354376
rect 176658 354320 176714 354356
rect 177578 352144 177634 352200
rect 176658 348064 176714 348120
rect 176658 345480 176714 345536
rect 176566 336504 176622 336560
rect 176474 332560 176530 332616
rect 176474 323584 176530 323640
rect 176658 334464 176714 334520
rect 176658 330384 176714 330440
rect 176658 325760 176714 325816
rect 177670 318824 177726 318880
rect 177578 316784 177634 316840
rect 176658 314880 176714 314936
rect 176658 312840 176714 312896
rect 176658 309984 176714 310040
rect 176658 303864 176714 303920
rect 176658 299240 176714 299296
rect 176658 297200 176714 297256
rect 176658 295160 176714 295216
rect 176658 290400 176714 290456
rect 176658 288380 176714 288416
rect 176658 288360 176660 288380
rect 176660 288360 176712 288380
rect 176712 288360 176714 288380
rect 176658 283600 176714 283656
rect 176658 281560 176714 281616
rect 176750 279520 176806 279576
rect 176658 277480 176714 277536
rect 176658 274760 176714 274816
rect 176658 272584 176714 272640
rect 176658 261840 176714 261896
rect 176658 256944 176714 257000
rect 176658 254904 176714 254960
rect 176658 252864 176714 252920
rect 176658 250824 176714 250880
rect 176658 246200 176714 246256
rect 177946 380296 178002 380352
rect 177946 309984 178002 310040
rect 177946 307944 178002 308000
rect 177854 305904 177910 305960
rect 177854 301144 177910 301200
rect 177762 270544 177818 270600
rect 179234 292304 179290 292360
rect 179142 263744 179198 263800
rect 178774 256672 178830 256728
rect 178774 226344 178830 226400
rect 190458 365744 190514 365800
rect 189998 360168 190054 360224
rect 179418 343304 179474 343360
rect 179326 286184 179382 286240
rect 179326 268504 179382 268560
rect 179510 341332 179566 341388
rect 208766 357584 208822 357640
rect 218058 378140 218114 378176
rect 218058 378120 218060 378140
rect 218060 378120 218112 378140
rect 218112 378120 218114 378140
rect 217046 358808 217102 358864
rect 222842 355272 222898 355328
rect 228822 356224 228878 356280
rect 233790 358944 233846 359000
rect 243266 532616 243322 532672
rect 244278 409128 244334 409184
rect 243542 407224 243598 407280
rect 245658 583208 245714 583264
rect 244554 515888 244610 515944
rect 245382 515888 245438 515944
rect 244554 445848 244610 445904
rect 245382 445848 245438 445904
rect 245290 409128 245346 409184
rect 245750 576408 245806 576464
rect 245750 573008 245806 573064
rect 245750 566208 245806 566264
rect 245750 560088 245806 560144
rect 245750 556688 245806 556744
rect 245750 549888 245806 549944
rect 245750 539688 245806 539744
rect 245934 569608 245990 569664
rect 245934 543088 245990 543144
rect 245842 536288 245898 536344
rect 245842 526088 245898 526144
rect 245842 522688 245898 522744
rect 245842 519288 245898 519344
rect 245842 512488 245898 512544
rect 245842 506404 245844 506424
rect 245844 506404 245896 506424
rect 245896 506404 245898 506424
rect 245842 506368 245898 506404
rect 245842 502968 245898 503024
rect 245842 499588 245898 499624
rect 245842 499568 245844 499588
rect 245844 499568 245896 499588
rect 245896 499568 245898 499588
rect 245842 496168 245898 496224
rect 245842 492768 245898 492824
rect 245842 485968 245898 486024
rect 245934 479168 245990 479224
rect 245842 475768 245898 475824
rect 245842 472368 245898 472424
rect 245934 462168 245990 462224
rect 245934 459448 245990 459504
rect 245934 456048 245990 456104
rect 246946 562808 247002 562864
rect 246670 509804 246672 509824
rect 246672 509804 246724 509824
rect 246724 509804 246726 509824
rect 246670 509768 246726 509804
rect 245934 449248 245990 449304
rect 246302 442448 246358 442504
rect 245934 439048 245990 439104
rect 245934 435648 245990 435704
rect 245934 432248 245990 432304
rect 245934 428848 245990 428904
rect 245934 425448 245990 425504
rect 245934 422048 245990 422104
rect 245934 418648 245990 418704
rect 245934 415248 245990 415304
rect 245934 411848 245990 411904
rect 246394 405728 246450 405784
rect 247130 482568 247186 482624
rect 244370 359352 244426 359408
rect 247222 465568 247278 465624
rect 249982 403688 250038 403744
rect 253938 583752 253994 583808
rect 253938 386960 253994 387016
rect 260838 586608 260894 586664
rect 254214 357584 254270 357640
rect 252466 356360 252522 356416
rect 263598 389952 263654 390008
rect 259458 367104 259514 367160
rect 260102 367104 260158 367160
rect 269762 367648 269818 367704
rect 292578 368872 292634 368928
rect 292578 368464 292634 368520
rect 291750 357448 291806 357504
rect 291290 354592 291346 354648
rect 292762 355952 292818 356008
rect 292394 354592 292450 354648
rect 293222 368872 293278 368928
rect 293130 355952 293186 356008
rect 293130 354728 293186 354784
rect 293038 350104 293094 350160
rect 293038 346976 293094 347032
rect 179510 262112 179566 262168
rect 179418 243616 179474 243672
rect 179602 244092 179658 244148
rect 179510 243480 179566 243536
rect 215298 240624 215354 240680
rect 179786 231784 179842 231840
rect 184202 237360 184258 237416
rect 194046 94832 194102 94888
rect 206282 177248 206338 177304
rect 213918 175616 213974 175672
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 213918 173576 213974 173632
rect 214010 172896 214066 172952
rect 213918 172216 213974 172272
rect 214102 171536 214158 171592
rect 213918 171028 213920 171048
rect 213920 171028 213972 171048
rect 213972 171028 213974 171048
rect 213918 170992 213974 171028
rect 214010 170312 214066 170368
rect 213918 168952 213974 169008
rect 214010 168292 214066 168328
rect 214010 168272 214012 168292
rect 214012 168272 214064 168292
rect 214064 168272 214066 168292
rect 213918 167592 213974 167648
rect 213918 166948 213920 166968
rect 213920 166948 213972 166968
rect 213972 166948 213974 166968
rect 213918 166912 213974 166948
rect 214010 166368 214066 166424
rect 213918 165688 213974 165744
rect 213918 165008 213974 165064
rect 214010 164328 214066 164384
rect 213918 162968 213974 163024
rect 213918 159704 213974 159760
rect 214010 159024 214066 159080
rect 213918 157664 213974 157720
rect 213918 157120 213974 157176
rect 214010 156440 214066 156496
rect 213918 155760 213974 155816
rect 214010 154400 214066 154456
rect 213918 153720 213974 153776
rect 214010 153040 214066 153096
rect 213918 152496 213974 152552
rect 214102 151136 214158 151192
rect 213918 150476 213974 150512
rect 213918 150456 213920 150476
rect 213920 150456 213972 150476
rect 213972 150456 213974 150476
rect 214010 149096 214066 149152
rect 213918 148416 213974 148472
rect 213918 147872 213974 147928
rect 213918 147192 213974 147248
rect 214654 161744 214710 161800
rect 214930 169632 214986 169688
rect 215022 161064 215078 161120
rect 214930 160384 214986 160440
rect 214654 151816 214710 151872
rect 214562 149776 214618 149832
rect 214562 146512 214618 146568
rect 213918 145832 213974 145888
rect 214470 145152 214526 145208
rect 213918 144472 213974 144528
rect 213918 143248 213974 143304
rect 213918 141888 213974 141944
rect 213182 141208 213238 141264
rect 214010 140528 214066 140584
rect 213918 139848 213974 139904
rect 214010 139168 214066 139224
rect 213918 138624 213974 138680
rect 214102 137944 214158 138000
rect 214930 142568 214986 142624
rect 214654 137264 214710 137320
rect 214010 136584 214066 136640
rect 213918 135904 213974 135960
rect 214562 135224 214618 135280
rect 213918 134544 213974 134600
rect 213918 132640 213974 132696
rect 214010 130600 214066 130656
rect 213918 129920 213974 129976
rect 213918 129240 213974 129296
rect 214010 128016 214066 128072
rect 213918 127336 213974 127392
rect 213918 126656 213974 126712
rect 214010 125296 214066 125352
rect 213918 124616 213974 124672
rect 214010 124072 214066 124128
rect 213918 123392 213974 123448
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 213274 121352 213330 121408
rect 213918 120672 213974 120728
rect 214102 119992 214158 120048
rect 214010 119448 214066 119504
rect 213918 118804 213920 118824
rect 213920 118804 213972 118824
rect 213972 118804 213974 118824
rect 213918 118768 213974 118804
rect 214010 118088 214066 118144
rect 213918 117408 213974 117464
rect 214010 116728 214066 116784
rect 213918 116048 213974 116104
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 214010 114144 214066 114200
rect 213918 113464 213974 113520
rect 214010 112784 214066 112840
rect 213918 112104 213974 112160
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 214010 110200 214066 110256
rect 213918 109520 213974 109576
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 214010 107480 214066 107536
rect 213918 106800 213974 106856
rect 214102 106120 214158 106176
rect 214010 105576 214066 105632
rect 213918 104932 213920 104952
rect 213920 104932 213972 104952
rect 213972 104932 213974 104952
rect 213918 104896 213974 104932
rect 214010 104216 214066 104272
rect 213918 103556 213974 103592
rect 213918 103536 213920 103556
rect 213920 103536 213972 103556
rect 213972 103536 213974 103556
rect 213918 102196 213974 102232
rect 213918 102176 213920 102196
rect 213920 102176 213972 102196
rect 213972 102176 213974 102196
rect 213918 100952 213974 101008
rect 214010 100272 214066 100328
rect 213918 99592 213974 99648
rect 214010 98912 214066 98968
rect 213918 98232 213974 98288
rect 213918 97552 213974 97608
rect 214838 131960 214894 132016
rect 214746 125976 214802 126032
rect 214746 102856 214802 102912
rect 214378 97144 214434 97200
rect 214654 96328 214710 96384
rect 214562 89120 214618 89176
rect 214930 101496 214986 101552
rect 214838 96872 214894 96928
rect 214746 89664 214802 89720
rect 224038 238720 224094 238776
rect 224958 191120 225014 191176
rect 229098 188536 229154 188592
rect 231122 178880 231178 178936
rect 239402 178744 239458 178800
rect 246394 177248 246450 177304
rect 248510 177520 248566 177576
rect 247682 176024 247738 176080
rect 248050 175752 248106 175808
rect 249154 175888 249210 175944
rect 249338 175208 249394 175264
rect 249154 174664 249210 174720
rect 249154 169088 249210 169144
rect 250442 186360 250498 186416
rect 249982 169496 250038 169552
rect 249890 149776 249946 149832
rect 249798 139440 249854 139496
rect 250534 136584 250590 136640
rect 252466 173712 252522 173768
rect 251730 172796 251732 172816
rect 251732 172796 251784 172816
rect 251784 172796 251786 172816
rect 251730 172760 251786 172796
rect 252466 172388 252468 172408
rect 252468 172388 252520 172408
rect 252520 172388 252522 172408
rect 252466 172352 252522 172388
rect 252558 171808 252614 171864
rect 252374 171400 252430 171456
rect 251546 170448 251602 170504
rect 252282 170040 252338 170096
rect 252190 168544 252246 168600
rect 252466 167592 252522 167648
rect 252282 167184 252338 167240
rect 252282 166640 252338 166696
rect 251914 166232 251970 166288
rect 252282 165688 252338 165744
rect 252466 165280 252522 165336
rect 251546 164328 251602 164384
rect 252466 163920 252522 163976
rect 252098 162968 252154 163024
rect 252466 162424 252522 162480
rect 252466 162016 252522 162072
rect 252466 161472 252522 161528
rect 252466 161084 252522 161120
rect 252466 161064 252468 161084
rect 252468 161064 252520 161084
rect 252520 161064 252522 161084
rect 252834 164192 252890 164248
rect 252742 160520 252798 160576
rect 252466 160112 252522 160168
rect 252466 159568 252522 159624
rect 251914 159160 251970 159216
rect 251454 158752 251510 158808
rect 252466 158208 252522 158264
rect 252466 157276 252522 157312
rect 252466 157256 252468 157276
rect 252468 157256 252520 157276
rect 252520 157256 252522 157276
rect 251546 156848 251602 156904
rect 251362 156304 251418 156360
rect 252466 155896 252522 155952
rect 251546 153992 251602 154048
rect 252374 154944 252430 155000
rect 252466 154420 252522 154456
rect 252466 154400 252468 154420
rect 252468 154400 252520 154420
rect 252520 154400 252522 154420
rect 252006 153448 252062 153504
rect 252466 153040 252522 153096
rect 252282 152632 252338 152688
rect 251730 152088 251786 152144
rect 251270 151136 251326 151192
rect 251270 146920 251326 146976
rect 251730 149232 251786 149288
rect 251546 148280 251602 148336
rect 251362 146512 251418 146568
rect 251730 146240 251786 146296
rect 251546 144064 251602 144120
rect 251730 143112 251786 143168
rect 251178 140800 251234 140856
rect 251178 140428 251180 140448
rect 251180 140428 251232 140448
rect 251232 140428 251234 140448
rect 251178 140392 251234 140428
rect 250810 137944 250866 138000
rect 251270 137536 251326 137592
rect 251730 135632 251786 135688
rect 251270 133320 251326 133376
rect 251730 131416 251786 131472
rect 252466 151680 252522 151736
rect 252374 150728 252430 150784
rect 252466 150184 252522 150240
rect 252466 148824 252522 148880
rect 252466 147464 252522 147520
rect 252466 145968 252522 146024
rect 252374 145560 252430 145616
rect 252098 145016 252154 145072
rect 252466 144608 252522 144664
rect 252098 143656 252154 143712
rect 251822 127200 251878 127256
rect 251730 126248 251786 126304
rect 251546 123936 251602 123992
rect 251270 122984 251326 123040
rect 251730 122032 251786 122088
rect 251730 120536 251786 120592
rect 251454 118768 251510 118824
rect 251730 117816 251786 117872
rect 251270 116864 251326 116920
rect 251546 115368 251602 115424
rect 251178 114960 251234 115016
rect 251730 112648 251786 112704
rect 251638 111152 251694 111208
rect 251546 110200 251602 110256
rect 252466 141752 252522 141808
rect 252374 141480 252430 141536
rect 252098 135224 252154 135280
rect 252282 134272 252338 134328
rect 251914 115912 251970 115968
rect 252834 141344 252890 141400
rect 252834 141072 252890 141128
rect 253202 139984 253258 140040
rect 252466 138488 252522 138544
rect 252466 136992 252522 137048
rect 252466 136176 252522 136232
rect 252466 134680 252522 134736
rect 252466 133764 252468 133784
rect 252468 133764 252520 133784
rect 252520 133764 252522 133784
rect 252466 133728 252522 133764
rect 252374 132776 252430 132832
rect 252190 132368 252246 132424
rect 252282 131824 252338 131880
rect 252466 130908 252468 130928
rect 252468 130908 252520 130928
rect 252520 130908 252522 130928
rect 252466 130872 252522 130908
rect 252374 130464 252430 130520
rect 252282 130056 252338 130112
rect 252466 129512 252522 129568
rect 252374 129104 252430 129160
rect 252282 128560 252338 128616
rect 252466 128188 252468 128208
rect 252468 128188 252520 128208
rect 252520 128188 252522 128208
rect 252466 128152 252522 128188
rect 252374 127608 252430 127664
rect 252466 126692 252468 126712
rect 252468 126692 252520 126712
rect 252520 126692 252522 126712
rect 252466 126656 252522 126692
rect 252190 125704 252246 125760
rect 252466 125296 252522 125352
rect 252098 124752 252154 124808
rect 252466 124344 252522 124400
rect 252466 123392 252522 123448
rect 252466 122440 252522 122496
rect 252374 121488 252430 121544
rect 252466 121080 252522 121136
rect 252374 120128 252430 120184
rect 252282 119584 252338 119640
rect 252190 119176 252246 119232
rect 252466 118224 252522 118280
rect 252282 117272 252338 117328
rect 252466 116320 252522 116376
rect 252466 114452 252468 114472
rect 252468 114452 252520 114472
rect 252520 114452 252522 114472
rect 252466 114416 252522 114452
rect 252374 114008 252430 114064
rect 252466 113464 252522 113520
rect 252098 112104 252154 112160
rect 252006 111696 252062 111752
rect 251822 106936 251878 106992
rect 251730 105032 251786 105088
rect 251178 102756 251180 102776
rect 251180 102756 251232 102776
rect 251232 102756 251234 102776
rect 251178 102720 251234 102756
rect 251178 101360 251234 101416
rect 251178 96600 251234 96656
rect 252098 110744 252154 110800
rect 252098 109248 252154 109304
rect 252190 108296 252246 108352
rect 252006 107888 252062 107944
rect 252098 106528 252154 106584
rect 252006 105984 252062 106040
rect 252190 104660 252192 104680
rect 252192 104660 252244 104680
rect 252244 104660 252246 104680
rect 252190 104624 252246 104660
rect 252466 109792 252522 109848
rect 252466 108876 252468 108896
rect 252468 108876 252520 108896
rect 252520 108876 252522 108896
rect 252466 108840 252522 108876
rect 252466 107500 252522 107536
rect 252466 107480 252468 107500
rect 252468 107480 252520 107500
rect 252520 107480 252522 107500
rect 252466 105576 252522 105632
rect 252374 104080 252430 104136
rect 252466 103672 252522 103728
rect 252282 103128 252338 103184
rect 252466 102176 252522 102232
rect 251914 101768 251970 101824
rect 251546 100408 251602 100464
rect 252006 99864 252062 99920
rect 251362 98912 251418 98968
rect 252466 100816 252522 100872
rect 252466 99456 252522 99512
rect 252466 98504 252522 98560
rect 254122 177248 254178 177304
rect 256790 169768 256846 169824
rect 252190 97008 252246 97064
rect 251362 96192 251418 96248
rect 261022 173848 261078 173904
rect 262218 222128 262274 222184
rect 262862 222128 262918 222184
rect 275282 235320 275338 235376
rect 269946 141344 270002 141400
rect 278318 3984 278374 4040
rect 283654 178608 283710 178664
rect 287702 240080 287758 240136
rect 292670 239148 292726 239184
rect 292670 239128 292672 239148
rect 292672 239128 292724 239148
rect 292724 239128 292726 239148
rect 293958 357312 294014 357368
rect 293314 354492 293316 354512
rect 293316 354492 293368 354512
rect 293368 354492 293370 354512
rect 293314 354456 293370 354492
rect 293958 352280 294014 352336
rect 293222 334600 293278 334656
rect 293130 314200 293186 314256
rect 293866 314200 293922 314256
rect 293130 287680 293186 287736
rect 293222 259120 293278 259176
rect 293314 241168 293370 241224
rect 294142 336640 294198 336696
rect 294050 331880 294106 331936
rect 294050 325760 294106 325816
rect 294142 312160 294198 312216
rect 295614 345480 295670 345536
rect 295614 340720 295670 340776
rect 295614 338680 295670 338736
rect 295522 327800 295578 327856
rect 295430 321000 295486 321056
rect 295430 318960 295486 319016
rect 295430 316920 295486 316976
rect 295338 310120 295394 310176
rect 294234 309032 294290 309088
rect 295522 308080 295578 308136
rect 295338 301280 295394 301336
rect 295338 299240 295394 299296
rect 295338 294480 295394 294536
rect 294234 267960 294290 268016
rect 295522 296520 295578 296576
rect 295614 292440 295670 292496
rect 295522 290400 295578 290456
rect 295430 285676 295432 285696
rect 295432 285676 295484 285696
rect 295484 285676 295486 285696
rect 295430 285640 295486 285676
rect 295430 283620 295486 283656
rect 295430 283600 295432 283620
rect 295432 283600 295484 283620
rect 295484 283600 295486 283620
rect 295430 281580 295486 281616
rect 295430 281560 295432 281580
rect 295432 281560 295484 281580
rect 295484 281560 295486 281580
rect 295430 278860 295486 278896
rect 295430 278840 295432 278860
rect 295432 278840 295484 278860
rect 295484 278840 295486 278860
rect 295430 276800 295486 276856
rect 295430 274760 295486 274816
rect 295430 272740 295486 272776
rect 295430 272720 295432 272740
rect 295432 272720 295484 272740
rect 295484 272720 295486 272740
rect 295430 270000 295486 270056
rect 295430 265920 295486 265976
rect 295522 263880 295578 263936
rect 295430 261160 295486 261216
rect 295522 255040 295578 255096
rect 295522 252320 295578 252376
rect 295522 250280 295578 250336
rect 295522 246200 295578 246256
rect 296626 343440 296682 343496
rect 296626 323040 296682 323096
rect 296902 329840 296958 329896
rect 296902 243480 296958 243536
rect 296074 3984 296130 4040
rect 301134 241032 301190 241088
rect 304262 354592 304318 354648
rect 307114 177248 307170 177304
rect 307022 175616 307078 175672
rect 307574 175208 307630 175264
rect 307022 174800 307078 174856
rect 306930 172216 306986 172272
rect 307298 174392 307354 174448
rect 307666 173984 307722 174040
rect 307574 173576 307630 173632
rect 307298 173168 307354 173224
rect 307666 172624 307722 172680
rect 307482 171808 307538 171864
rect 307390 170992 307446 171048
rect 307298 169804 307300 169824
rect 307300 169804 307352 169824
rect 307352 169804 307354 169824
rect 307298 169768 307354 169804
rect 307298 168428 307354 168464
rect 307298 168408 307300 168428
rect 307300 168408 307352 168428
rect 307352 168408 307354 168428
rect 307114 168000 307170 168056
rect 306930 167592 306986 167648
rect 306930 166776 306986 166832
rect 305642 162832 305698 162888
rect 307022 161608 307078 161664
rect 306746 161200 306802 161256
rect 306930 158616 306986 158672
rect 306746 156984 306802 157040
rect 306654 153176 306710 153232
rect 306562 152224 306618 152280
rect 306930 150184 306986 150240
rect 306746 147192 306802 147248
rect 307482 170584 307538 170640
rect 307666 170176 307722 170232
rect 307574 169224 307630 169280
rect 307666 168816 307722 168872
rect 307206 167184 307262 167240
rect 307666 166368 307722 166424
rect 307482 165824 307538 165880
rect 307574 165416 307630 165472
rect 307390 165008 307446 165064
rect 307298 164228 307300 164248
rect 307300 164228 307352 164248
rect 307352 164228 307354 164248
rect 307298 164192 307354 164228
rect 307298 163376 307354 163432
rect 307666 164600 307722 164656
rect 307574 163784 307630 163840
rect 307666 162968 307722 163024
rect 307574 162832 307630 162888
rect 307482 162424 307538 162480
rect 307666 162016 307722 162072
rect 307482 160792 307538 160848
rect 307666 160384 307722 160440
rect 307574 159976 307630 160032
rect 307206 159024 307262 159080
rect 307666 159568 307722 159624
rect 307666 158208 307722 158264
rect 307298 157800 307354 157856
rect 307666 157392 307722 157448
rect 307482 156576 307538 156632
rect 307390 156168 307446 156224
rect 307482 155624 307538 155680
rect 307574 155216 307630 155272
rect 307666 154808 307722 154864
rect 307482 154400 307538 154456
rect 307666 153992 307722 154048
rect 307574 153584 307630 153640
rect 307482 152632 307538 152688
rect 307666 151836 307722 151872
rect 307666 151816 307668 151836
rect 307668 151816 307720 151836
rect 307720 151816 307722 151836
rect 307482 151408 307538 151464
rect 307390 150592 307446 150648
rect 307298 149252 307354 149288
rect 307298 149232 307300 149252
rect 307300 149232 307352 149252
rect 307352 149232 307354 149252
rect 307114 148008 307170 148064
rect 306930 144608 306986 144664
rect 306562 144200 306618 144256
rect 306746 142976 306802 143032
rect 307022 141208 307078 141264
rect 306930 136584 306986 136640
rect 305734 134408 305790 134464
rect 305642 124616 305698 124672
rect 304354 115096 304410 115152
rect 306930 133592 306986 133648
rect 306562 133184 306618 133240
rect 306930 132232 306986 132288
rect 306746 129240 306802 129296
rect 306562 126384 306618 126440
rect 306930 125840 306986 125896
rect 306930 125432 306986 125488
rect 306930 121624 306986 121680
rect 306746 121216 306802 121272
rect 306930 119992 306986 120048
rect 306562 119584 306618 119640
rect 307298 147600 307354 147656
rect 307206 145424 307262 145480
rect 307114 130600 307170 130656
rect 306562 118224 306618 118280
rect 306746 117000 306802 117056
rect 306746 115640 306802 115696
rect 307022 114008 307078 114064
rect 306930 108024 306986 108080
rect 305826 107752 305882 107808
rect 305918 105168 305974 105224
rect 306746 103400 306802 103456
rect 306562 101632 306618 101688
rect 306746 97824 306802 97880
rect 307298 142432 307354 142488
rect 307666 151000 307722 151056
rect 307482 149776 307538 149832
rect 307666 148824 307722 148880
rect 307482 148416 307538 148472
rect 307666 146784 307722 146840
rect 307574 146376 307630 146432
rect 307482 145832 307538 145888
rect 307666 145016 307722 145072
rect 307482 143792 307538 143848
rect 307666 143384 307722 143440
rect 307574 142024 307630 142080
rect 307482 141616 307538 141672
rect 307666 140800 307722 140856
rect 307666 139576 307722 139632
rect 307482 139032 307538 139088
rect 307574 138624 307630 138680
rect 307666 138216 307722 138272
rect 307574 137808 307630 137864
rect 307482 137400 307538 137456
rect 307666 136992 307722 137048
rect 307482 136176 307538 136232
rect 307666 135632 307722 135688
rect 307482 134816 307538 134872
rect 307666 134020 307722 134056
rect 307666 134000 307668 134020
rect 307668 134000 307720 134020
rect 307720 134000 307722 134020
rect 307666 132660 307722 132696
rect 307666 132640 307668 132660
rect 307668 132640 307720 132660
rect 307720 132640 307722 132660
rect 307666 131824 307722 131880
rect 307390 131416 307446 131472
rect 307298 129820 307300 129840
rect 307300 129820 307352 129840
rect 307352 129820 307354 129840
rect 307298 129784 307354 129820
rect 307298 128444 307354 128480
rect 307298 128424 307300 128444
rect 307300 128424 307352 128444
rect 307352 128424 307354 128444
rect 307666 130192 307722 130248
rect 307666 128832 307722 128888
rect 307574 127608 307630 127664
rect 307666 127200 307722 127256
rect 307482 125024 307538 125080
rect 307666 124244 307668 124264
rect 307668 124244 307720 124264
rect 307720 124244 307722 124264
rect 307666 124208 307722 124244
rect 307574 123800 307630 123856
rect 307482 122984 307538 123040
rect 307666 123392 307722 123448
rect 307206 96192 307262 96248
rect 307482 122440 307538 122496
rect 307666 122032 307722 122088
rect 307482 120808 307538 120864
rect 307666 120400 307722 120456
rect 307666 119040 307722 119096
rect 307574 118632 307630 118688
rect 307666 117816 307722 117872
rect 307574 116592 307630 116648
rect 307666 116184 307722 116240
rect 307574 115232 307630 115288
rect 307666 114824 307722 114880
rect 307574 113600 307630 113656
rect 307666 113228 307668 113248
rect 307668 113228 307720 113248
rect 307720 113228 307722 113248
rect 307666 113192 307722 113228
rect 307482 112648 307538 112704
rect 307574 112240 307630 112296
rect 307666 111832 307722 111888
rect 307482 111424 307538 111480
rect 307666 111016 307722 111072
rect 307574 110608 307630 110664
rect 307482 110200 307538 110256
rect 307574 109792 307630 109848
rect 307666 109248 307722 109304
rect 307482 108840 307538 108896
rect 307574 108432 307630 108488
rect 307482 107752 307538 107808
rect 307666 107616 307722 107672
rect 307482 107208 307538 107264
rect 307574 106800 307630 106856
rect 307666 106392 307722 106448
rect 307666 105848 307722 105904
rect 307482 105440 307538 105496
rect 307666 105168 307722 105224
rect 307666 105032 307722 105088
rect 307574 104624 307630 104680
rect 307482 104216 307538 104272
rect 307666 103808 307722 103864
rect 307482 102992 307538 103048
rect 307666 102448 307722 102504
rect 308218 102040 308274 102096
rect 308218 101088 308274 101144
rect 307666 100816 307722 100872
rect 307574 100408 307630 100464
rect 307666 99592 307722 99648
rect 307666 99048 307722 99104
rect 307574 98640 307630 98696
rect 307482 98232 307538 98288
rect 307482 97416 307538 97472
rect 307666 96600 307722 96656
rect 301962 6160 302018 6216
rect 303158 3440 303214 3496
rect 307942 3440 307998 3496
rect 308678 139984 308734 140040
rect 308678 139440 308734 139496
rect 309046 3984 309102 4040
rect 314658 238720 314714 238776
rect 314566 235184 314622 235240
rect 318154 177384 318210 177440
rect 323030 235184 323086 235240
rect 318430 176568 318486 176624
rect 318246 176160 318302 176216
rect 321466 176024 321522 176080
rect 321282 170312 321338 170368
rect 321742 174392 321798 174448
rect 321834 172624 321890 172680
rect 321650 148280 321706 148336
rect 321650 107480 321706 107536
rect 321558 105984 321614 106040
rect 321558 102176 321614 102232
rect 321374 97280 321430 97336
rect 321374 95920 321430 95976
rect 321466 95804 321522 95840
rect 321466 95784 321468 95804
rect 321468 95784 321520 95804
rect 321520 95784 321522 95804
rect 310518 79328 310574 79384
rect 323030 176568 323086 176624
rect 323030 173168 323086 173224
rect 324318 223624 324374 223680
rect 324410 193840 324466 193896
rect 324318 170892 324320 170912
rect 324320 170892 324372 170912
rect 324372 170892 324374 170912
rect 324318 170856 324374 170892
rect 324318 168544 324374 168600
rect 324502 174664 324558 174720
rect 324410 167728 324466 167784
rect 324318 167048 324374 167104
rect 324318 165452 324320 165472
rect 324320 165452 324372 165472
rect 324372 165452 324374 165472
rect 324318 165416 324374 165452
rect 324410 164736 324466 164792
rect 324318 163920 324374 163976
rect 324410 163104 324466 163160
rect 324318 161608 324374 161664
rect 324318 160112 324374 160168
rect 324318 159296 324374 159352
rect 324318 158480 324374 158536
rect 324410 157800 324466 157856
rect 324318 156984 324374 157040
rect 324410 156304 324466 156360
rect 324962 223624 325018 223680
rect 325698 210296 325754 210352
rect 324594 155488 324650 155544
rect 324318 154672 324374 154728
rect 324318 153992 324374 154048
rect 324410 153176 324466 153232
rect 324318 152360 324374 152416
rect 324318 151700 324374 151736
rect 324318 151680 324320 151700
rect 324320 151680 324372 151700
rect 324372 151680 324374 151700
rect 324410 150864 324466 150920
rect 324318 149368 324374 149424
rect 324318 148552 324374 148608
rect 324318 147056 324374 147112
rect 323674 146240 323730 146296
rect 324318 144744 324374 144800
rect 324318 143112 324374 143168
rect 324318 138488 324374 138544
rect 324318 137808 324374 137864
rect 324318 134680 324374 134736
rect 324318 133184 324374 133240
rect 324502 136992 324558 137048
rect 324502 134000 324558 134056
rect 324318 132404 324320 132424
rect 324320 132404 324372 132424
rect 324372 132404 324374 132424
rect 324318 132368 324374 132404
rect 324410 131688 324466 131744
rect 324410 130872 324466 130928
rect 324318 130056 324374 130112
rect 324318 129376 324374 129432
rect 324410 128560 324466 128616
rect 324318 127744 324374 127800
rect 324410 127064 324466 127120
rect 324318 126248 324374 126304
rect 324502 125432 324558 125488
rect 325606 124752 325662 124808
rect 327078 219272 327134 219328
rect 325790 145424 325846 145480
rect 325974 177520 326030 177576
rect 325882 136312 325938 136368
rect 324318 123120 324374 123176
rect 324318 122440 324374 122496
rect 324410 121624 324466 121680
rect 324318 120808 324374 120864
rect 328550 227704 328606 227760
rect 329838 220768 329894 220824
rect 327170 142024 327226 142080
rect 324410 120128 324466 120184
rect 324318 119312 324374 119368
rect 324318 118532 324320 118552
rect 324320 118532 324372 118552
rect 324372 118532 324374 118552
rect 324318 118496 324374 118532
rect 324410 117816 324466 117872
rect 323490 116456 323546 116512
rect 323490 115912 323546 115968
rect 324318 115504 324374 115560
rect 324410 114688 324466 114744
rect 324318 114008 324374 114064
rect 324410 113192 324466 113248
rect 324318 112376 324374 112432
rect 324318 111732 324320 111752
rect 324320 111732 324372 111752
rect 324372 111732 324374 111752
rect 324318 111696 324374 111732
rect 324410 110880 324466 110936
rect 324318 110064 324374 110120
rect 323122 108568 323178 108624
rect 323030 107072 323086 107128
rect 322938 106256 322994 106312
rect 321742 104216 321798 104272
rect 322938 100816 322994 100872
rect 321834 98096 321890 98152
rect 310242 3304 310298 3360
rect 324318 103944 324374 104000
rect 324318 103128 324374 103184
rect 324318 101632 324374 101688
rect 324502 100136 324558 100192
rect 324410 99320 324466 99376
rect 324594 97008 324650 97064
rect 324410 93744 324466 93800
rect 324594 92384 324650 92440
rect 319718 3576 319774 3632
rect 331310 88984 331366 89040
rect 332690 21256 332746 21312
rect 336738 221992 336794 222048
rect 336738 196696 336794 196752
rect 336922 184184 336978 184240
rect 339498 202136 339554 202192
rect 339682 188264 339738 188320
rect 339866 1944 339922 2000
rect 342166 3440 342222 3496
rect 342442 200640 342498 200696
rect 342626 179152 342682 179208
rect 343914 179968 343970 180024
rect 346306 179324 346308 179344
rect 346308 179324 346360 179344
rect 346360 179324 346362 179344
rect 346306 179288 346362 179324
rect 345662 18672 345718 18728
rect 347778 50224 347834 50280
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580262 617480 580318 617536
rect 580170 590960 580226 591016
rect 579802 577632 579858 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580354 524456 580410 524512
rect 580078 471416 580134 471472
rect 580170 458088 580226 458144
rect 580170 418240 580226 418296
rect 582378 431568 582434 431624
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 395342 375264 395398 375320
rect 580906 365064 580962 365120
rect 580262 351872 580318 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 258848 580226 258904
rect 580170 245520 580226 245576
rect 580262 240760 580318 240816
rect 580170 232328 580226 232384
rect 580170 219000 580226 219056
rect 579894 205672 579950 205728
rect 580354 226888 580410 226944
rect 580354 192480 580410 192536
rect 580262 179152 580318 179208
rect 582562 354456 582618 354512
rect 582470 272176 582526 272232
rect 582470 238584 582526 238640
rect 582378 152632 582434 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 579618 39208 579674 39264
rect 579894 33108 579950 33144
rect 579894 33088 579896 33108
rect 579896 33088 579948 33108
rect 579948 33088 579950 33108
rect 579894 19760 579950 19816
rect 582562 165824 582618 165880
rect 582470 6568 582526 6624
<< obsm2 >>
rect 68800 95100 164756 174600
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580257 617538 580323 617541
rect 583520 617538 584960 617628
rect 580257 617536 584960 617538
rect 580257 617480 580262 617536
rect 580318 617480 584960 617536
rect 580257 617478 584960 617480
rect 580257 617475 580323 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect 58617 586666 58683 586669
rect 83365 586666 83431 586669
rect 58617 586664 83431 586666
rect 58617 586608 58622 586664
rect 58678 586608 83370 586664
rect 83426 586608 83431 586664
rect 58617 586606 83431 586608
rect 58617 586603 58683 586606
rect 83365 586603 83431 586606
rect 232773 586666 232839 586669
rect 260833 586666 260899 586669
rect 232773 586664 260899 586666
rect 232773 586608 232778 586664
rect 232834 586608 260838 586664
rect 260894 586608 260899 586664
rect 232773 586606 260899 586608
rect 232773 586603 232839 586606
rect 260833 586603 260899 586606
rect 243486 586468 243492 586532
rect 243556 586468 243562 586532
rect 41321 586394 41387 586397
rect 99373 586394 99439 586397
rect 41321 586392 99439 586394
rect 41321 586336 41326 586392
rect 41382 586336 99378 586392
rect 99434 586336 99439 586392
rect 41321 586334 99439 586336
rect 41321 586331 41387 586334
rect 99373 586331 99439 586334
rect 201401 586394 201467 586397
rect 243494 586394 243554 586468
rect 201401 586392 243554 586394
rect 201401 586336 201406 586392
rect 201462 586336 243554 586392
rect 201401 586334 243554 586336
rect 201401 586331 201467 586334
rect 169661 585442 169727 585445
rect 247166 585442 247172 585444
rect 169661 585440 247172 585442
rect 169661 585384 169666 585440
rect 169722 585384 247172 585440
rect 169661 585382 247172 585384
rect 169661 585379 169727 585382
rect 247166 585380 247172 585382
rect 247236 585380 247242 585444
rect 50981 585306 51047 585309
rect 178677 585306 178743 585309
rect 50981 585304 178743 585306
rect 50981 585248 50986 585304
rect 51042 585248 178682 585304
rect 178738 585248 178743 585304
rect 50981 585246 178743 585248
rect 50981 585243 51047 585246
rect 178677 585243 178743 585246
rect 61377 585170 61443 585173
rect 243261 585170 243327 585173
rect 61377 585168 243327 585170
rect 61377 585112 61382 585168
rect 61438 585112 243266 585168
rect 243322 585112 243327 585168
rect 61377 585110 243327 585112
rect 61377 585107 61443 585110
rect 243261 585107 243327 585110
rect 243629 585172 243695 585173
rect 243629 585168 243676 585172
rect 243740 585170 243746 585172
rect 243629 585112 243634 585168
rect 243629 585108 243676 585112
rect 243740 585110 243786 585170
rect 243740 585108 243746 585110
rect 243629 585107 243695 585108
rect 63534 584564 63540 584628
rect 63604 584626 63610 584628
rect 64413 584626 64479 584629
rect 92749 584626 92815 584629
rect 188061 584626 188127 584629
rect 63604 584624 64479 584626
rect 63604 584568 64418 584624
rect 64474 584568 64479 584624
rect 63604 584566 64479 584568
rect 63604 584564 63610 584566
rect 64413 584563 64479 584566
rect 84150 584624 92815 584626
rect 84150 584568 92754 584624
rect 92810 584568 92815 584624
rect 84150 584566 92815 584568
rect 50838 583884 50844 583948
rect 50908 583946 50914 583948
rect 84150 583946 84210 584566
rect 92749 584563 92815 584566
rect 180750 584624 188127 584626
rect 180750 584568 188066 584624
rect 188122 584568 188127 584624
rect 180750 584566 188127 584568
rect 50908 583886 84210 583946
rect 50908 583884 50914 583886
rect 57789 583810 57855 583813
rect 180750 583810 180810 584566
rect 188061 584563 188127 584566
rect 223481 584626 223547 584629
rect 223481 584624 229110 584626
rect 223481 584568 223486 584624
rect 223542 584568 229110 584624
rect 223481 584566 229110 584568
rect 223481 584563 223547 584566
rect 57789 583808 180810 583810
rect 57789 583752 57794 583808
rect 57850 583752 180810 583808
rect 57789 583750 180810 583752
rect 229050 583810 229110 584566
rect 253933 583810 253999 583813
rect 229050 583808 253999 583810
rect 229050 583752 253938 583808
rect 253994 583752 253999 583808
rect 229050 583750 253999 583752
rect 57789 583747 57855 583750
rect 253933 583747 253999 583750
rect 245653 583266 245719 583269
rect 243892 583264 245719 583266
rect 243892 583208 245658 583264
rect 245714 583208 245719 583264
rect 243892 583206 245719 583208
rect 245653 583203 245719 583206
rect 58934 582524 58940 582588
rect 59004 582586 59010 582588
rect 59004 582526 64124 582586
rect 59004 582524 59010 582526
rect 243537 580954 243603 580957
rect 243670 580954 243676 580956
rect 243537 580952 243676 580954
rect 243537 580896 243542 580952
rect 243598 580896 243676 580952
rect 243537 580894 243676 580896
rect 243537 580891 243603 580894
rect 243670 580892 243676 580894
rect 243740 580892 243746 580956
rect -960 580002 480 580092
rect 2865 580002 2931 580005
rect -960 580000 2931 580002
rect -960 579944 2870 580000
rect 2926 579944 2931 580000
rect -960 579942 2931 579944
rect -960 579852 480 579942
rect 2865 579939 2931 579942
rect 243310 579596 243370 579836
rect 243302 579532 243308 579596
rect 243372 579532 243378 579596
rect 57830 579124 57836 579188
rect 57900 579186 57906 579188
rect 57900 579126 64124 579186
rect 57900 579124 57906 579126
rect 243486 578852 243492 578916
rect 243556 578914 243562 578916
rect 295374 578914 295380 578916
rect 243556 578854 295380 578914
rect 243556 578852 243562 578854
rect 295374 578852 295380 578854
rect 295444 578852 295450 578916
rect 579797 577690 579863 577693
rect 583520 577690 584960 577780
rect 579797 577688 584960 577690
rect 579797 577632 579802 577688
rect 579858 577632 584960 577688
rect 579797 577630 584960 577632
rect 579797 577627 579863 577630
rect 583520 577540 584960 577630
rect 245745 576466 245811 576469
rect 243892 576464 245811 576466
rect 243892 576408 245750 576464
rect 245806 576408 245811 576464
rect 243892 576406 245811 576408
rect 245745 576403 245811 576406
rect 60038 575724 60044 575788
rect 60108 575786 60114 575788
rect 60108 575726 64124 575786
rect 60108 575724 60114 575726
rect 245745 573066 245811 573069
rect 243892 573064 245811 573066
rect 243892 573008 245750 573064
rect 245806 573008 245811 573064
rect 243892 573006 245811 573008
rect 245745 573003 245811 573006
rect 61878 572324 61884 572388
rect 61948 572386 61954 572388
rect 61948 572326 64124 572386
rect 61948 572324 61954 572326
rect 245929 569666 245995 569669
rect 246982 569666 246988 569668
rect 243892 569664 246988 569666
rect 243892 569608 245934 569664
rect 245990 569608 246988 569664
rect 243892 569606 246988 569608
rect 245929 569603 245995 569606
rect 246982 569604 246988 569606
rect 247052 569604 247058 569668
rect 60733 568986 60799 568989
rect 60733 568984 64124 568986
rect 60733 568928 60738 568984
rect 60794 568928 64124 568984
rect 60733 568926 64124 568928
rect 60733 568923 60799 568926
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 245745 566266 245811 566269
rect 243892 566264 245811 566266
rect 243892 566208 245750 566264
rect 245806 566208 245811 566264
rect 243892 566206 245811 566208
rect 245745 566203 245811 566206
rect 60733 565586 60799 565589
rect 60733 565584 64124 565586
rect 60733 565528 60738 565584
rect 60794 565528 64124 565584
rect 60733 565526 64124 565528
rect 60733 565523 60799 565526
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 246941 562866 247007 562869
rect 243892 562864 247007 562866
rect 243892 562808 246946 562864
rect 247002 562808 247007 562864
rect 243892 562806 247007 562808
rect 246941 562803 247007 562806
rect 60733 562186 60799 562189
rect 60733 562184 64124 562186
rect 60733 562128 60738 562184
rect 60794 562128 64124 562184
rect 60733 562126 64124 562128
rect 60733 562123 60799 562126
rect 245745 560146 245811 560149
rect 243892 560144 245811 560146
rect 243892 560088 245750 560144
rect 245806 560088 245811 560144
rect 243892 560086 245811 560088
rect 245745 560083 245811 560086
rect 31661 558242 31727 558245
rect 63534 558242 63540 558244
rect 31661 558240 63540 558242
rect 31661 558184 31666 558240
rect 31722 558184 63540 558240
rect 31661 558182 63540 558184
rect 31661 558179 31727 558182
rect 63534 558180 63540 558182
rect 63604 558180 63610 558244
rect 54334 557500 54340 557564
rect 54404 557562 54410 557564
rect 64094 557562 64154 558756
rect 54404 557502 64154 557562
rect 54404 557500 54410 557502
rect 245745 556746 245811 556749
rect 243892 556744 245811 556746
rect 243892 556688 245750 556744
rect 245806 556688 245811 556744
rect 243892 556686 245811 556688
rect 245745 556683 245811 556686
rect 60733 555386 60799 555389
rect 60733 555384 64124 555386
rect 60733 555328 60738 555384
rect 60794 555328 64124 555384
rect 60733 555326 64124 555328
rect 60733 555323 60799 555326
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 244222 553346 244228 553348
rect 243892 553286 244228 553346
rect 244222 553284 244228 553286
rect 244292 553284 244298 553348
rect 60733 552666 60799 552669
rect 60733 552664 64124 552666
rect 60733 552608 60738 552664
rect 60794 552608 64124 552664
rect 60733 552606 64124 552608
rect 60733 552603 60799 552606
rect 583520 551020 584960 551260
rect 245745 549946 245811 549949
rect 243892 549944 245811 549946
rect 243892 549888 245750 549944
rect 245806 549888 245811 549944
rect 243892 549886 245811 549888
rect 245745 549883 245811 549886
rect 60733 549266 60799 549269
rect 60733 549264 64124 549266
rect 60733 549208 60738 549264
rect 60794 549208 64124 549264
rect 60733 549206 64124 549208
rect 60733 549203 60799 549206
rect 244406 546546 244412 546548
rect 243892 546486 244412 546546
rect 244406 546484 244412 546486
rect 244476 546484 244482 546548
rect 62021 545866 62087 545869
rect 62021 545864 64124 545866
rect 62021 545808 62026 545864
rect 62082 545808 64124 545864
rect 62021 545806 64124 545808
rect 62021 545803 62087 545806
rect 245929 543146 245995 543149
rect 243892 543144 245995 543146
rect 243892 543088 245934 543144
rect 245990 543088 245995 543144
rect 243892 543086 245995 543088
rect 245929 543083 245995 543086
rect 60733 542466 60799 542469
rect 60733 542464 64124 542466
rect 60733 542408 60738 542464
rect 60794 542408 64124 542464
rect 60733 542406 64124 542408
rect 60733 542403 60799 542406
rect -960 540684 480 540924
rect 245745 539746 245811 539749
rect 243892 539744 245811 539746
rect 243892 539688 245750 539744
rect 245806 539688 245811 539744
rect 243892 539686 245811 539688
rect 245745 539683 245811 539686
rect 60733 539066 60799 539069
rect 60733 539064 64124 539066
rect 60733 539008 60738 539064
rect 60794 539008 64124 539064
rect 60733 539006 64124 539008
rect 60733 539003 60799 539006
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect 245837 536346 245903 536349
rect 243892 536344 245903 536346
rect 243892 536288 245842 536344
rect 245898 536288 245903 536344
rect 243892 536286 245903 536288
rect 245837 536283 245903 536286
rect 60733 535666 60799 535669
rect 60733 535664 64124 535666
rect 60733 535608 60738 535664
rect 60794 535608 64124 535664
rect 60733 535606 64124 535608
rect 60733 535603 60799 535606
rect 243310 532677 243370 532916
rect 243261 532672 243370 532677
rect 243261 532616 243266 532672
rect 243322 532616 243370 532672
rect 243261 532614 243370 532616
rect 243261 532611 243327 532614
rect 55622 532204 55628 532268
rect 55692 532266 55698 532268
rect 55692 532206 64124 532266
rect 55692 532204 55698 532206
rect 245694 529546 245700 529548
rect 243892 529486 245700 529546
rect 245694 529484 245700 529486
rect 245764 529484 245770 529548
rect 60733 528866 60799 528869
rect 60733 528864 64124 528866
rect 60733 528808 60738 528864
rect 60794 528808 64124 528864
rect 60733 528806 64124 528808
rect 60733 528803 60799 528806
rect -960 527914 480 528004
rect 3693 527914 3759 527917
rect -960 527912 3759 527914
rect -960 527856 3698 527912
rect 3754 527856 3759 527912
rect -960 527854 3759 527856
rect -960 527764 480 527854
rect 3693 527851 3759 527854
rect 245837 526146 245903 526149
rect 243892 526144 245903 526146
rect 243892 526088 245842 526144
rect 245898 526088 245903 526144
rect 243892 526086 245903 526088
rect 245837 526083 245903 526086
rect 59118 525404 59124 525468
rect 59188 525466 59194 525468
rect 63309 525466 63375 525469
rect 59188 525464 64124 525466
rect 59188 525408 63314 525464
rect 63370 525408 64124 525464
rect 59188 525406 64124 525408
rect 59188 525404 59194 525406
rect 63309 525403 63375 525406
rect 580349 524514 580415 524517
rect 583520 524514 584960 524604
rect 580349 524512 584960 524514
rect 580349 524456 580354 524512
rect 580410 524456 584960 524512
rect 580349 524454 584960 524456
rect 580349 524451 580415 524454
rect 583520 524364 584960 524454
rect 245837 522746 245903 522749
rect 243892 522744 245903 522746
rect 243892 522688 245842 522744
rect 245898 522688 245903 522744
rect 243892 522686 245903 522688
rect 245837 522683 245903 522686
rect 61653 522066 61719 522069
rect 61653 522064 64124 522066
rect 61653 522008 61658 522064
rect 61714 522008 64124 522064
rect 61653 522006 64124 522008
rect 61653 522003 61719 522006
rect 245837 519346 245903 519349
rect 243892 519344 245903 519346
rect 243892 519288 245842 519344
rect 245898 519288 245903 519344
rect 243892 519286 245903 519288
rect 245837 519283 245903 519286
rect 60365 518666 60431 518669
rect 60365 518664 64124 518666
rect 60365 518608 60370 518664
rect 60426 518608 64124 518664
rect 60365 518606 64124 518608
rect 60365 518603 60431 518606
rect 244549 515946 244615 515949
rect 245377 515946 245443 515949
rect 243892 515944 245443 515946
rect 243892 515888 244554 515944
rect 244610 515888 245382 515944
rect 245438 515888 245443 515944
rect 243892 515886 245443 515888
rect 244549 515883 244615 515886
rect 245377 515883 245443 515886
rect 60733 515266 60799 515269
rect 60733 515264 64124 515266
rect 60733 515208 60738 515264
rect 60794 515208 64124 515264
rect 60733 515206 64124 515208
rect 60733 515203 60799 515206
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 245837 512546 245903 512549
rect 243892 512544 245903 512546
rect 243892 512488 245842 512544
rect 245898 512488 245903 512544
rect 243892 512486 245903 512488
rect 245837 512483 245903 512486
rect 63534 511804 63540 511868
rect 63604 511866 63610 511868
rect 63604 511806 64124 511866
rect 63604 511804 63610 511806
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 61929 510506 61995 510509
rect 62062 510506 62068 510508
rect 61929 510504 62068 510506
rect 61929 510448 61934 510504
rect 61990 510448 62068 510504
rect 61929 510446 62068 510448
rect 61929 510443 61995 510446
rect 62062 510444 62068 510446
rect 62132 510444 62138 510508
rect 246665 509826 246731 509829
rect 243892 509824 246731 509826
rect 243892 509768 246670 509824
rect 246726 509768 246731 509824
rect 243892 509766 246731 509768
rect 246665 509763 246731 509766
rect 61929 508466 61995 508469
rect 61929 508464 64124 508466
rect 61929 508408 61934 508464
rect 61990 508408 64124 508464
rect 61929 508406 64124 508408
rect 61929 508403 61995 508406
rect 245837 506426 245903 506429
rect 243892 506424 245903 506426
rect 243892 506368 245842 506424
rect 245898 506368 245903 506424
rect 243892 506366 245903 506368
rect 245837 506363 245903 506366
rect 60549 505066 60615 505069
rect 60549 505064 64124 505066
rect 60549 505008 60554 505064
rect 60610 505008 64124 505064
rect 60549 505006 64124 505008
rect 60549 505003 60615 505006
rect 245837 503026 245903 503029
rect 243892 503024 245903 503026
rect 243892 502968 245842 503024
rect 245898 502968 245903 503024
rect 243892 502966 245903 502968
rect 245837 502963 245903 502966
rect 60733 502346 60799 502349
rect 60733 502344 64124 502346
rect 60733 502288 60738 502344
rect 60794 502288 64124 502344
rect 60733 502286 64124 502288
rect 60733 502283 60799 502286
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 245837 499626 245903 499629
rect 243892 499624 245903 499626
rect 243892 499568 245842 499624
rect 245898 499568 245903 499624
rect 243892 499566 245903 499568
rect 245837 499563 245903 499566
rect 63033 498946 63099 498949
rect 63033 498944 64124 498946
rect 63033 498888 63038 498944
rect 63094 498888 64124 498944
rect 63033 498886 64124 498888
rect 63033 498883 63099 498886
rect 583520 497844 584960 498084
rect 245837 496226 245903 496229
rect 243892 496224 245903 496226
rect 243892 496168 245842 496224
rect 245898 496168 245903 496224
rect 243892 496166 245903 496168
rect 245837 496163 245903 496166
rect 60733 495546 60799 495549
rect 60733 495544 64124 495546
rect 60733 495488 60738 495544
rect 60794 495488 64124 495544
rect 60733 495486 64124 495488
rect 60733 495483 60799 495486
rect 245837 492826 245903 492829
rect 243892 492824 245903 492826
rect 243892 492768 245842 492824
rect 245898 492768 245903 492824
rect 243892 492766 245903 492768
rect 245837 492763 245903 492766
rect 60733 492146 60799 492149
rect 60733 492144 64124 492146
rect 60733 492088 60738 492144
rect 60794 492088 64124 492144
rect 60733 492086 64124 492088
rect 60733 492083 60799 492086
rect 245878 489426 245884 489428
rect 243892 489366 245884 489426
rect 245878 489364 245884 489366
rect 245948 489364 245954 489428
rect -960 488596 480 488836
rect 60733 488746 60799 488749
rect 60733 488744 64124 488746
rect 60733 488688 60738 488744
rect 60794 488688 64124 488744
rect 60733 488686 64124 488688
rect 60733 488683 60799 488686
rect 245837 486026 245903 486029
rect 243892 486024 245903 486026
rect 243892 485968 245842 486024
rect 245898 485968 245903 486024
rect 243892 485966 245903 485968
rect 245837 485963 245903 485966
rect 61837 485890 61903 485893
rect 62062 485890 62068 485892
rect 61837 485888 62068 485890
rect 61837 485832 61842 485888
rect 61898 485832 62068 485888
rect 61837 485830 62068 485832
rect 61837 485827 61903 485830
rect 62062 485828 62068 485830
rect 62132 485828 62138 485892
rect 61193 485346 61259 485349
rect 61193 485344 64124 485346
rect 61193 485288 61198 485344
rect 61254 485288 64124 485344
rect 61193 485286 64124 485288
rect 61193 485283 61259 485286
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 247125 482626 247191 482629
rect 243892 482624 247191 482626
rect 243892 482568 247130 482624
rect 247186 482568 247191 482624
rect 243892 482566 247191 482568
rect 247125 482563 247191 482566
rect 61561 481946 61627 481949
rect 61561 481944 64124 481946
rect 61561 481888 61566 481944
rect 61622 481888 64124 481944
rect 61561 481886 64124 481888
rect 61561 481883 61627 481886
rect 245929 479226 245995 479229
rect 243892 479224 245995 479226
rect 243892 479168 245934 479224
rect 245990 479168 245995 479224
rect 243892 479166 245995 479168
rect 245929 479163 245995 479166
rect 60733 478546 60799 478549
rect 60733 478544 64124 478546
rect 60733 478488 60738 478544
rect 60794 478488 64124 478544
rect 60733 478486 64124 478488
rect 60733 478483 60799 478486
rect 245837 475826 245903 475829
rect 243892 475824 245903 475826
rect -960 475690 480 475780
rect 243892 475768 245842 475824
rect 245898 475768 245903 475824
rect 243892 475766 245903 475768
rect 245837 475763 245903 475766
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 61377 475146 61443 475149
rect 61377 475144 64124 475146
rect 61377 475088 61382 475144
rect 61438 475088 64124 475144
rect 61377 475086 64124 475088
rect 61377 475083 61443 475086
rect 61837 473242 61903 473245
rect 63718 473242 63724 473244
rect 61837 473240 63724 473242
rect 61837 473184 61842 473240
rect 61898 473184 63724 473240
rect 61837 473182 63724 473184
rect 61837 473179 61903 473182
rect 63718 473180 63724 473182
rect 63788 473180 63794 473244
rect 245837 472426 245903 472429
rect 243892 472424 245903 472426
rect 243892 472368 245842 472424
rect 245898 472368 245903 472424
rect 243892 472366 245903 472368
rect 245837 472363 245903 472366
rect 60917 471746 60983 471749
rect 63493 471746 63559 471749
rect 60917 471744 64124 471746
rect 60917 471688 60922 471744
rect 60978 471688 63498 471744
rect 63554 471688 64124 471744
rect 60917 471686 64124 471688
rect 60917 471683 60983 471686
rect 63493 471683 63559 471686
rect 580073 471474 580139 471477
rect 583520 471474 584960 471564
rect 580073 471472 584960 471474
rect 580073 471416 580078 471472
rect 580134 471416 584960 471472
rect 580073 471414 584960 471416
rect 580073 471411 580139 471414
rect 583520 471324 584960 471414
rect 49550 469780 49556 469844
rect 49620 469842 49626 469844
rect 58617 469842 58683 469845
rect 49620 469840 58683 469842
rect 49620 469784 58622 469840
rect 58678 469784 58683 469840
rect 49620 469782 58683 469784
rect 49620 469780 49626 469782
rect 58617 469779 58683 469782
rect 60733 468346 60799 468349
rect 243862 468346 243922 468996
rect 60733 468344 64124 468346
rect 60733 468288 60738 468344
rect 60794 468288 64124 468344
rect 60733 468286 64124 468288
rect 243862 468286 248430 468346
rect 60733 468283 60799 468286
rect 248370 467938 248430 468286
rect 328494 467938 328500 467940
rect 248370 467878 328500 467938
rect 328494 467876 328500 467878
rect 328564 467876 328570 467940
rect 247217 465626 247283 465629
rect 243892 465624 247283 465626
rect 243892 465568 247222 465624
rect 247278 465568 247283 465624
rect 243892 465566 247283 465568
rect 247217 465563 247283 465566
rect 53598 464884 53604 464948
rect 53668 464946 53674 464948
rect 53741 464946 53807 464949
rect 53668 464944 53807 464946
rect 53668 464888 53746 464944
rect 53802 464888 53807 464944
rect 53668 464886 53807 464888
rect 53668 464884 53674 464886
rect 53741 464883 53807 464886
rect 60733 464946 60799 464949
rect 60733 464944 64124 464946
rect 60733 464888 60738 464944
rect 60794 464888 64124 464944
rect 60733 464886 64124 464888
rect 60733 464883 60799 464886
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 245929 462226 245995 462229
rect 243892 462224 245995 462226
rect 243892 462168 245934 462224
rect 245990 462168 245995 462224
rect 243892 462166 245995 462168
rect 245929 462163 245995 462166
rect 60733 461546 60799 461549
rect 60733 461544 64124 461546
rect 60733 461488 60738 461544
rect 60794 461488 64124 461544
rect 60733 461486 64124 461488
rect 60733 461483 60799 461486
rect 245929 459506 245995 459509
rect 243892 459504 245995 459506
rect 243892 459448 245934 459504
rect 245990 459448 245995 459504
rect 243892 459446 245995 459448
rect 245929 459443 245995 459446
rect 60733 458146 60799 458149
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 60733 458144 64124 458146
rect 60733 458088 60738 458144
rect 60794 458088 64124 458144
rect 60733 458086 64124 458088
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 60733 458083 60799 458086
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 245929 456106 245995 456109
rect 243892 456104 245995 456106
rect 243892 456048 245934 456104
rect 245990 456048 245995 456104
rect 243892 456046 245995 456048
rect 245929 456043 245995 456046
rect 61745 454746 61811 454749
rect 61745 454744 64124 454746
rect 61745 454688 61750 454744
rect 61806 454688 64124 454744
rect 61745 454686 64124 454688
rect 61745 454683 61811 454686
rect 331254 452706 331260 452708
rect 243892 452646 331260 452706
rect 331254 452644 331260 452646
rect 331324 452644 331330 452708
rect 61837 452026 61903 452029
rect 61837 452024 64124 452026
rect 61837 451968 61842 452024
rect 61898 451968 64124 452024
rect 61837 451966 64124 451968
rect 61837 451963 61903 451966
rect 63309 449986 63375 449989
rect 63718 449986 63724 449988
rect 63309 449984 63724 449986
rect 63309 449928 63314 449984
rect 63370 449928 63724 449984
rect 63309 449926 63724 449928
rect 63309 449923 63375 449926
rect 63718 449924 63724 449926
rect 63788 449924 63794 449988
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 245929 449306 245995 449309
rect 243892 449304 245995 449306
rect 243892 449248 245934 449304
rect 245990 449248 245995 449304
rect 243892 449246 245995 449248
rect 245929 449243 245995 449246
rect 63350 448564 63356 448628
rect 63420 448626 63426 448628
rect 63420 448566 64124 448626
rect 63420 448564 63426 448566
rect 244549 445906 244615 445909
rect 245377 445906 245443 445909
rect 243892 445904 245443 445906
rect 243892 445848 244554 445904
rect 244610 445848 245382 445904
rect 245438 445848 245443 445904
rect 243892 445846 245443 445848
rect 244549 445843 244615 445846
rect 245377 445843 245443 445846
rect 60733 445226 60799 445229
rect 60733 445224 64124 445226
rect 60733 445168 60738 445224
rect 60794 445168 64124 445224
rect 60733 445166 64124 445168
rect 60733 445163 60799 445166
rect 583520 444668 584960 444908
rect 246297 442506 246363 442509
rect 243892 442504 246363 442506
rect 243892 442448 246302 442504
rect 246358 442448 246363 442504
rect 243892 442446 246363 442448
rect 246297 442443 246363 442446
rect 60733 441826 60799 441829
rect 60733 441824 64124 441826
rect 60733 441768 60738 441824
rect 60794 441768 64124 441824
rect 60733 441766 64124 441768
rect 60733 441763 60799 441766
rect 245929 439106 245995 439109
rect 243892 439104 245995 439106
rect 243892 439048 245934 439104
rect 245990 439048 245995 439104
rect 243892 439046 245995 439048
rect 245929 439043 245995 439046
rect 60917 438426 60983 438429
rect 63401 438426 63467 438429
rect 60917 438424 64124 438426
rect 60917 438368 60922 438424
rect 60978 438368 63406 438424
rect 63462 438368 64124 438424
rect 60917 438366 64124 438368
rect 60917 438363 60983 438366
rect 63401 438363 63467 438366
rect -960 436508 480 436748
rect 245929 435706 245995 435709
rect 243892 435704 245995 435706
rect 243892 435648 245934 435704
rect 245990 435648 245995 435704
rect 243892 435646 245995 435648
rect 245929 435643 245995 435646
rect 61561 435026 61627 435029
rect 61561 435024 64124 435026
rect 61561 434968 61566 435024
rect 61622 434968 64124 435024
rect 61561 434966 64124 434968
rect 61561 434963 61627 434966
rect 57646 434556 57652 434620
rect 57716 434618 57722 434620
rect 58709 434618 58775 434621
rect 57716 434616 58775 434618
rect 57716 434560 58714 434616
rect 58770 434560 58775 434616
rect 57716 434558 58775 434560
rect 57716 434556 57722 434558
rect 58709 434555 58775 434558
rect 245929 432306 245995 432309
rect 243892 432304 245995 432306
rect 243892 432248 245934 432304
rect 245990 432248 245995 432304
rect 243892 432246 245995 432248
rect 245929 432243 245995 432246
rect 582373 431626 582439 431629
rect 583520 431626 584960 431716
rect 582373 431624 584960 431626
rect 53414 430612 53420 430676
rect 53484 430674 53490 430676
rect 64094 430674 64154 431596
rect 582373 431568 582378 431624
rect 582434 431568 584960 431624
rect 582373 431566 584960 431568
rect 582373 431563 582439 431566
rect 583520 431476 584960 431566
rect 53484 430614 64154 430674
rect 53484 430612 53490 430614
rect 63217 429314 63283 429317
rect 64086 429314 64092 429316
rect 63217 429312 64092 429314
rect 63217 429256 63222 429312
rect 63278 429256 64092 429312
rect 63217 429254 64092 429256
rect 63217 429251 63283 429254
rect 64086 429252 64092 429254
rect 64156 429252 64162 429316
rect 245929 428906 245995 428909
rect 243892 428904 245995 428906
rect 243892 428848 245934 428904
rect 245990 428848 245995 428904
rect 243892 428846 245995 428848
rect 245929 428843 245995 428846
rect 60733 428226 60799 428229
rect 60733 428224 64124 428226
rect 60733 428168 60738 428224
rect 60794 428168 64124 428224
rect 60733 428166 64124 428168
rect 60733 428163 60799 428166
rect 245929 425506 245995 425509
rect 243892 425504 245995 425506
rect 243892 425448 245934 425504
rect 245990 425448 245995 425504
rect 243892 425446 245995 425448
rect 245929 425443 245995 425446
rect 60733 424826 60799 424829
rect 60733 424824 64124 424826
rect 60733 424768 60738 424824
rect 60794 424768 64124 424824
rect 60733 424766 64124 424768
rect 60733 424763 60799 424766
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 245929 422106 245995 422109
rect 243892 422104 245995 422106
rect 243892 422048 245934 422104
rect 245990 422048 245995 422104
rect 243892 422046 245995 422048
rect 245929 422043 245995 422046
rect 63166 421364 63172 421428
rect 63236 421426 63242 421428
rect 63236 421366 64124 421426
rect 63236 421364 63242 421366
rect 245929 418706 245995 418709
rect 243892 418704 245995 418706
rect 243892 418648 245934 418704
rect 245990 418648 245995 418704
rect 243892 418646 245995 418648
rect 245929 418643 245995 418646
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 62297 418026 62363 418029
rect 62297 418024 64124 418026
rect 62297 417968 62302 418024
rect 62358 417968 64124 418024
rect 62297 417966 64124 417968
rect 62297 417963 62363 417966
rect 245929 415306 245995 415309
rect 243892 415304 245995 415306
rect 243892 415248 245934 415304
rect 245990 415248 245995 415304
rect 243892 415246 245995 415248
rect 245929 415243 245995 415246
rect 60733 414626 60799 414629
rect 60733 414624 64124 414626
rect 60733 414568 60738 414624
rect 60794 414568 64124 414624
rect 60733 414566 64124 414568
rect 60733 414563 60799 414566
rect 245929 411906 245995 411909
rect 243892 411904 245995 411906
rect 243892 411848 245934 411904
rect 245990 411848 245995 411904
rect 243892 411846 245995 411848
rect 245929 411843 245995 411846
rect 63677 410682 63743 410685
rect 64094 410682 64154 411196
rect 63677 410680 64154 410682
rect -960 410546 480 410636
rect 63677 410624 63682 410680
rect 63738 410624 64154 410680
rect 63677 410622 64154 410624
rect 63677 410619 63743 410622
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 244273 409186 244339 409189
rect 245285 409186 245351 409189
rect 243892 409184 245351 409186
rect 243892 409128 244278 409184
rect 244334 409128 245290 409184
rect 245346 409128 245351 409184
rect 243892 409126 245351 409128
rect 244273 409123 244339 409126
rect 245285 409123 245351 409126
rect 60733 407826 60799 407829
rect 60733 407824 64124 407826
rect 60733 407768 60738 407824
rect 60794 407768 64124 407824
rect 60733 407766 64124 407768
rect 60733 407763 60799 407766
rect 243302 407220 243308 407284
rect 243372 407282 243378 407284
rect 243537 407282 243603 407285
rect 243372 407280 243603 407282
rect 243372 407224 243542 407280
rect 243598 407224 243603 407280
rect 243372 407222 243603 407224
rect 243372 407220 243378 407222
rect 243537 407219 243603 407222
rect 246389 405786 246455 405789
rect 243892 405784 246455 405786
rect 243892 405728 246394 405784
rect 246450 405728 246455 405784
rect 243892 405726 246455 405728
rect 246389 405723 246455 405726
rect 53414 405588 53420 405652
rect 53484 405650 53490 405652
rect 53557 405650 53623 405653
rect 53484 405648 53623 405650
rect 53484 405592 53562 405648
rect 53618 405592 53623 405648
rect 53484 405590 53623 405592
rect 53484 405588 53490 405590
rect 53557 405587 53623 405590
rect 242801 405514 242867 405517
rect 247166 405514 247172 405516
rect 242801 405512 247172 405514
rect 242801 405456 242806 405512
rect 242862 405456 247172 405512
rect 242801 405454 247172 405456
rect 242801 405451 242867 405454
rect 247166 405452 247172 405454
rect 247236 405452 247242 405516
rect 57646 404908 57652 404972
rect 57716 404970 57722 404972
rect 73153 404970 73219 404973
rect 57716 404968 73219 404970
rect 57716 404912 73158 404968
rect 73214 404912 73219 404968
rect 57716 404910 73219 404912
rect 57716 404908 57722 404910
rect 73153 404907 73219 404910
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 63166 404500 63172 404564
rect 63236 404562 63242 404564
rect 66161 404562 66227 404565
rect 63236 404560 66227 404562
rect 63236 404504 66166 404560
rect 66222 404504 66227 404560
rect 63236 404502 66227 404504
rect 63236 404500 63242 404502
rect 66161 404499 66227 404502
rect 61878 404364 61884 404428
rect 61948 404426 61954 404428
rect 65517 404426 65583 404429
rect 61948 404424 65583 404426
rect 61948 404368 65522 404424
rect 65578 404368 65583 404424
rect 61948 404366 65583 404368
rect 61948 404364 61954 404366
rect 65517 404363 65583 404366
rect 44081 403746 44147 403749
rect 66846 403746 66852 403748
rect 44081 403744 66852 403746
rect 44081 403688 44086 403744
rect 44142 403688 66852 403744
rect 44081 403686 66852 403688
rect 44081 403683 44147 403686
rect 66846 403684 66852 403686
rect 66916 403684 66922 403748
rect 176561 403746 176627 403749
rect 249977 403746 250043 403749
rect 176561 403744 250043 403746
rect 176561 403688 176566 403744
rect 176622 403688 249982 403744
rect 250038 403688 250043 403744
rect 176561 403686 250043 403688
rect 176561 403683 176627 403686
rect 249977 403683 250043 403686
rect 54937 403610 55003 403613
rect 103513 403610 103579 403613
rect 54937 403608 103579 403610
rect 54937 403552 54942 403608
rect 54998 403552 103518 403608
rect 103574 403552 103579 403608
rect 54937 403550 103579 403552
rect 54937 403547 55003 403550
rect 103513 403547 103579 403550
rect 159357 403610 159423 403613
rect 243302 403610 243308 403612
rect 159357 403608 243308 403610
rect 159357 403552 159362 403608
rect 159418 403552 243308 403608
rect 159357 403550 243308 403552
rect 159357 403547 159423 403550
rect 243302 403548 243308 403550
rect 243372 403548 243378 403612
rect 52361 401706 52427 401709
rect 52494 401706 52500 401708
rect 52361 401704 52500 401706
rect 52361 401648 52366 401704
rect 52422 401648 52500 401704
rect 52361 401646 52500 401648
rect 52361 401643 52427 401646
rect 52494 401644 52500 401646
rect 52564 401644 52570 401708
rect 147581 401026 147647 401029
rect 245878 401026 245884 401028
rect 147581 401024 245884 401026
rect 147581 400968 147586 401024
rect 147642 400968 245884 401024
rect 147581 400966 245884 400968
rect 147581 400963 147647 400966
rect 245878 400964 245884 400966
rect 245948 400964 245954 401028
rect 118601 400890 118667 400893
rect 244406 400890 244412 400892
rect 118601 400888 244412 400890
rect 118601 400832 118606 400888
rect 118662 400832 244412 400888
rect 118601 400830 244412 400832
rect 118601 400827 118667 400830
rect 244406 400828 244412 400830
rect 244476 400828 244482 400892
rect 58934 399468 58940 399532
rect 59004 399530 59010 399532
rect 67633 399530 67699 399533
rect 59004 399528 67699 399530
rect 59004 399472 67638 399528
rect 67694 399472 67699 399528
rect 59004 399470 67699 399472
rect 59004 399468 59010 399470
rect 67633 399467 67699 399470
rect 50838 398108 50844 398172
rect 50908 398170 50914 398172
rect 76005 398170 76071 398173
rect 50908 398168 76071 398170
rect 50908 398112 76010 398168
rect 76066 398112 76071 398168
rect 50908 398110 76071 398112
rect 50908 398108 50914 398110
rect 76005 398107 76071 398110
rect 63534 397972 63540 398036
rect 63604 398034 63610 398036
rect 90357 398034 90423 398037
rect 63604 398032 90423 398034
rect 63604 397976 90362 398032
rect 90418 397976 90423 398032
rect 63604 397974 90423 397976
rect 63604 397972 63610 397974
rect 90357 397971 90423 397974
rect -960 397490 480 397580
rect 3969 397490 4035 397493
rect -960 397488 4035 397490
rect -960 397432 3974 397488
rect 4030 397432 4035 397488
rect -960 397430 4035 397432
rect -960 397340 480 397430
rect 3969 397427 4035 397430
rect 583520 391628 584960 391868
rect 180006 389948 180012 390012
rect 180076 390010 180082 390012
rect 263593 390010 263659 390013
rect 180076 390008 263659 390010
rect 180076 389952 263598 390008
rect 263654 389952 263659 390008
rect 180076 389950 263659 389952
rect 180076 389948 180082 389950
rect 263593 389947 263659 389950
rect 108941 389874 109007 389877
rect 244222 389874 244228 389876
rect 108941 389872 244228 389874
rect 108941 389816 108946 389872
rect 109002 389816 244228 389872
rect 108941 389814 244228 389816
rect 108941 389811 109007 389814
rect 244222 389812 244228 389814
rect 244292 389812 244298 389876
rect 60038 386956 60044 387020
rect 60108 387018 60114 387020
rect 105537 387018 105603 387021
rect 60108 387016 105603 387018
rect 60108 386960 105542 387016
rect 105598 386960 105603 387016
rect 60108 386958 105603 386960
rect 60108 386956 60114 386958
rect 105537 386955 105603 386958
rect 178534 386956 178540 387020
rect 178604 387018 178610 387020
rect 253933 387018 253999 387021
rect 178604 387016 253999 387018
rect 178604 386960 253938 387016
rect 253994 386960 253999 387016
rect 178604 386958 253999 386960
rect 178604 386956 178610 386958
rect 253933 386955 253999 386958
rect -960 384284 480 384524
rect 177941 380354 178007 380357
rect 246982 380354 246988 380356
rect 177941 380352 246988 380354
rect 177941 380296 177946 380352
rect 178002 380296 246988 380352
rect 177941 380294 246988 380296
rect 177941 380291 178007 380294
rect 246982 380292 246988 380294
rect 247052 380292 247058 380356
rect 95877 380218 95943 380221
rect 242934 380218 242940 380220
rect 95877 380216 242940 380218
rect 95877 380160 95882 380216
rect 95938 380160 242940 380216
rect 95877 380158 242940 380160
rect 95877 380155 95943 380158
rect 242934 380156 242940 380158
rect 243004 380156 243010 380220
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 70894 378116 70900 378180
rect 70964 378178 70970 378180
rect 218053 378178 218119 378181
rect 70964 378176 218119 378178
rect 70964 378120 218058 378176
rect 218114 378120 218119 378176
rect 70964 378118 218119 378120
rect 70964 378116 70970 378118
rect 218053 378115 218119 378118
rect 151813 376682 151879 376685
rect 152549 376682 152615 376685
rect 151813 376680 152615 376682
rect 151813 376624 151818 376680
rect 151874 376624 152554 376680
rect 152610 376624 152615 376680
rect 151813 376622 152615 376624
rect 151813 376619 151879 376622
rect 152549 376619 152615 376622
rect 152549 375458 152615 375461
rect 152549 375456 293970 375458
rect 152549 375400 152554 375456
rect 152610 375400 293970 375456
rect 152549 375398 293970 375400
rect 152549 375395 152615 375398
rect 293910 375322 293970 375398
rect 295006 375322 295012 375324
rect 293910 375262 295012 375322
rect 295006 375260 295012 375262
rect 295076 375322 295082 375324
rect 395337 375322 395403 375325
rect 295076 375320 395403 375322
rect 295076 375264 395342 375320
rect 395398 375264 395403 375320
rect 295076 375262 395403 375264
rect 295076 375260 295082 375262
rect 395337 375259 395403 375262
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 292573 368930 292639 368933
rect 293217 368930 293283 368933
rect 292573 368928 293283 368930
rect 292573 368872 292578 368928
rect 292634 368872 293222 368928
rect 293278 368872 293283 368928
rect 292573 368870 293283 368872
rect 292573 368867 292639 368870
rect 293217 368867 293283 368870
rect 146886 368460 146892 368524
rect 146956 368522 146962 368524
rect 292573 368522 292639 368525
rect 146956 368520 292639 368522
rect 146956 368464 292578 368520
rect 292634 368464 292639 368520
rect 146956 368462 292639 368464
rect 146956 368460 146962 368462
rect 292573 368459 292639 368462
rect 269757 367706 269823 367709
rect 295558 367706 295564 367708
rect 269757 367704 295564 367706
rect 269757 367648 269762 367704
rect 269818 367648 295564 367704
rect 269757 367646 295564 367648
rect 269757 367643 269823 367646
rect 295558 367644 295564 367646
rect 295628 367644 295634 367708
rect 134374 367100 134380 367164
rect 134444 367162 134450 367164
rect 259453 367162 259519 367165
rect 260097 367162 260163 367165
rect 134444 367160 260163 367162
rect 134444 367104 259458 367160
rect 259514 367104 260102 367160
rect 260158 367104 260163 367160
rect 134444 367102 260163 367104
rect 134444 367100 134450 367102
rect 259453 367099 259519 367102
rect 260097 367099 260163 367102
rect 190453 365802 190519 365805
rect 332542 365802 332548 365804
rect 190453 365800 332548 365802
rect 190453 365744 190458 365800
rect 190514 365744 332548 365800
rect 190453 365742 332548 365744
rect 190453 365739 190519 365742
rect 332542 365740 332548 365742
rect 332612 365740 332618 365804
rect 580901 365122 580967 365125
rect 583520 365122 584960 365212
rect 580901 365120 584960 365122
rect 580901 365064 580906 365120
rect 580962 365064 584960 365120
rect 580901 365062 584960 365064
rect 580901 365059 580967 365062
rect 583520 364972 584960 365062
rect 131021 362266 131087 362269
rect 245694 362266 245700 362268
rect 131021 362264 245700 362266
rect 131021 362208 131026 362264
rect 131082 362208 245700 362264
rect 131021 362206 245700 362208
rect 131021 362203 131087 362206
rect 245694 362204 245700 362206
rect 245764 362204 245770 362268
rect 189993 360226 190059 360229
rect 340822 360226 340828 360228
rect 189993 360224 340828 360226
rect 189993 360168 189998 360224
rect 190054 360168 340828 360224
rect 189993 360166 340828 360168
rect 189993 360163 190059 360166
rect 340822 360164 340828 360166
rect 340892 360164 340898 360228
rect 61837 359410 61903 359413
rect 119654 359410 119660 359412
rect 61837 359408 119660 359410
rect 61837 359352 61842 359408
rect 61898 359352 119660 359408
rect 61837 359350 119660 359352
rect 61837 359347 61903 359350
rect 119654 359348 119660 359350
rect 119724 359348 119730 359412
rect 172278 359348 172284 359412
rect 172348 359410 172354 359412
rect 244365 359410 244431 359413
rect 172348 359408 244431 359410
rect 172348 359352 244370 359408
rect 244426 359352 244431 359408
rect 172348 359350 244431 359352
rect 172348 359348 172354 359350
rect 244365 359347 244431 359350
rect 233785 359002 233851 359005
rect 299974 359002 299980 359004
rect 233785 359000 299980 359002
rect 233785 358944 233790 359000
rect 233846 358944 299980 359000
rect 233785 358942 299980 358944
rect 233785 358939 233851 358942
rect 299974 358940 299980 358942
rect 300044 358940 300050 359004
rect 217041 358866 217107 358869
rect 296478 358866 296484 358868
rect 217041 358864 296484 358866
rect 217041 358808 217046 358864
rect 217102 358808 296484 358864
rect 217041 358806 296484 358808
rect 217041 358803 217107 358806
rect 296478 358804 296484 358806
rect 296548 358804 296554 358868
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 39849 358050 39915 358053
rect 161749 358050 161815 358053
rect 39849 358048 161815 358050
rect 39849 357992 39854 358048
rect 39910 357992 161754 358048
rect 161810 357992 161815 358048
rect 39849 357990 161815 357992
rect 39849 357987 39915 357990
rect 161749 357987 161815 357990
rect 129038 357580 129044 357644
rect 129108 357642 129114 357644
rect 208761 357642 208827 357645
rect 129108 357640 208827 357642
rect 129108 357584 208766 357640
rect 208822 357584 208827 357640
rect 129108 357582 208827 357584
rect 129108 357580 129114 357582
rect 208761 357579 208827 357582
rect 254209 357642 254275 357645
rect 298502 357642 298508 357644
rect 254209 357640 298508 357642
rect 254209 357584 254214 357640
rect 254270 357584 298508 357640
rect 254209 357582 298508 357584
rect 254209 357579 254275 357582
rect 298502 357580 298508 357582
rect 298572 357580 298578 357644
rect 161473 357506 161539 357509
rect 161749 357506 161815 357509
rect 291745 357506 291811 357509
rect 161473 357504 291811 357506
rect 161473 357448 161478 357504
rect 161534 357448 161754 357504
rect 161810 357448 291750 357504
rect 291806 357448 291811 357504
rect 161473 357446 291811 357448
rect 161473 357443 161539 357446
rect 161749 357443 161815 357446
rect 291745 357443 291811 357446
rect 293953 357372 294019 357373
rect 293902 357370 293908 357372
rect 293862 357310 293908 357370
rect 293972 357368 294019 357372
rect 294014 357312 294019 357368
rect 293902 357308 293908 357310
rect 293972 357308 294019 357312
rect 293953 357307 294019 357308
rect 64086 356628 64092 356692
rect 64156 356690 64162 356692
rect 64156 356630 122850 356690
rect 64156 356628 64162 356630
rect 122790 356146 122850 356630
rect 252461 356418 252527 356421
rect 301446 356418 301452 356420
rect 252461 356416 301452 356418
rect 252461 356360 252466 356416
rect 252522 356360 301452 356416
rect 252461 356358 301452 356360
rect 252461 356355 252527 356358
rect 301446 356356 301452 356358
rect 301516 356356 301522 356420
rect 228817 356282 228883 356285
rect 304206 356282 304212 356284
rect 228817 356280 304212 356282
rect 228817 356224 228822 356280
rect 228878 356224 304212 356280
rect 228817 356222 304212 356224
rect 228817 356219 228883 356222
rect 304206 356220 304212 356222
rect 304276 356220 304282 356284
rect 132585 356146 132651 356149
rect 292614 356146 292620 356148
rect 122790 356144 292620 356146
rect 122790 356088 132590 356144
rect 132646 356088 292620 356144
rect 122790 356086 292620 356088
rect 132585 356083 132651 356086
rect 292614 356084 292620 356086
rect 292684 356084 292690 356148
rect 292757 356010 292823 356013
rect 293125 356010 293191 356013
rect 292757 356008 293191 356010
rect 292757 355952 292762 356008
rect 292818 355952 293130 356008
rect 293186 355952 293191 356008
rect 292757 355950 293191 355952
rect 292757 355947 292823 355950
rect 293125 355947 293191 355950
rect 177062 355268 177068 355332
rect 177132 355330 177138 355332
rect 222837 355330 222903 355333
rect 177132 355328 222903 355330
rect 177132 355272 222842 355328
rect 222898 355272 222903 355328
rect 177132 355270 222903 355272
rect 177132 355268 177138 355270
rect 222837 355267 222903 355270
rect 113173 354786 113239 354789
rect 293125 354786 293191 354789
rect 113173 354784 293191 354786
rect 113173 354728 113178 354784
rect 113234 354728 293130 354784
rect 293186 354728 293191 354784
rect 113173 354726 293191 354728
rect 113173 354723 113239 354726
rect 293125 354723 293191 354726
rect 53598 354588 53604 354652
rect 53668 354650 53674 354652
rect 165429 354650 165495 354653
rect 53668 354648 165495 354650
rect 53668 354592 165434 354648
rect 165490 354592 165495 354648
rect 53668 354590 165495 354592
rect 53668 354588 53674 354590
rect 165429 354587 165495 354590
rect 291285 354650 291351 354653
rect 292389 354650 292455 354653
rect 304257 354650 304323 354653
rect 291285 354648 292314 354650
rect 291285 354592 291290 354648
rect 291346 354592 292314 354648
rect 291285 354590 292314 354592
rect 291285 354587 291351 354590
rect 176653 354378 176719 354381
rect 176653 354376 180044 354378
rect 176653 354320 176658 354376
rect 176714 354320 180044 354376
rect 292254 354348 292314 354590
rect 292389 354648 304323 354650
rect 292389 354592 292394 354648
rect 292450 354592 304262 354648
rect 304318 354592 304323 354648
rect 292389 354590 304323 354592
rect 292389 354587 292455 354590
rect 304257 354587 304323 354590
rect 293309 354514 293375 354517
rect 582557 354514 582623 354517
rect 293309 354512 582623 354514
rect 293309 354456 293314 354512
rect 293370 354456 582562 354512
rect 582618 354456 582623 354512
rect 293309 354454 582623 354456
rect 293309 354451 293375 354454
rect 582557 354451 582623 354454
rect 176653 354318 180044 354320
rect 176653 354315 176719 354318
rect 164233 353426 164299 353429
rect 165429 353426 165495 353429
rect 164233 353424 165495 353426
rect 164233 353368 164238 353424
rect 164294 353368 165434 353424
rect 165490 353368 165495 353424
rect 164233 353366 165495 353368
rect 164233 353363 164299 353366
rect 165429 353363 165495 353366
rect 152406 352548 152412 352612
rect 152476 352610 152482 352612
rect 179822 352610 179828 352612
rect 152476 352550 179828 352610
rect 152476 352548 152482 352550
rect 179822 352548 179828 352550
rect 179892 352548 179898 352612
rect 293953 352338 294019 352341
rect 292836 352336 294019 352338
rect 292836 352280 293958 352336
rect 294014 352280 294019 352336
rect 292836 352278 294019 352280
rect 293953 352275 294019 352278
rect 179462 352210 180044 352270
rect 177573 352202 177639 352205
rect 179462 352202 179522 352210
rect 177573 352200 179522 352202
rect 177573 352144 177578 352200
rect 177634 352144 179522 352200
rect 177573 352142 179522 352144
rect 177573 352139 177639 352142
rect 580257 351930 580323 351933
rect 583520 351930 584960 352020
rect 580257 351928 584960 351930
rect 580257 351872 580262 351928
rect 580318 351872 584960 351928
rect 580257 351870 584960 351872
rect 580257 351867 580323 351870
rect 583520 351780 584960 351870
rect 179462 350170 180044 350230
rect 176510 350100 176516 350164
rect 176580 350162 176586 350164
rect 179462 350162 179522 350170
rect 293033 350162 293099 350165
rect 176580 350102 179522 350162
rect 292806 350160 293099 350162
rect 292806 350104 293038 350160
rect 293094 350104 293099 350160
rect 292806 350102 293099 350104
rect 176580 350100 176586 350102
rect 110321 349754 110387 349757
rect 178534 349754 178540 349756
rect 110321 349752 178540 349754
rect 110321 349696 110326 349752
rect 110382 349696 178540 349752
rect 110321 349694 178540 349696
rect 110321 349691 110387 349694
rect 178534 349692 178540 349694
rect 178604 349692 178610 349756
rect 292806 349588 292866 350102
rect 293033 350099 293099 350102
rect 179462 348130 180044 348190
rect 176653 348122 176719 348125
rect 179462 348122 179522 348130
rect 176653 348120 179522 348122
rect 176653 348064 176658 348120
rect 176714 348064 179522 348120
rect 176653 348062 179522 348064
rect 176653 348059 176719 348062
rect 292806 347034 292866 347548
rect 293033 347034 293099 347037
rect 292806 347032 293099 347034
rect 292806 346976 293038 347032
rect 293094 346976 293099 347032
rect 292806 346974 293099 346976
rect 293033 346971 293099 346974
rect 176653 345538 176719 345541
rect 295609 345538 295675 345541
rect 176653 345536 179522 345538
rect -960 345402 480 345492
rect 176653 345480 176658 345536
rect 176714 345480 179522 345536
rect 176653 345478 179522 345480
rect 292836 345536 295675 345538
rect 292836 345480 295614 345536
rect 295670 345480 295675 345536
rect 292836 345478 295675 345480
rect 176653 345475 176719 345478
rect 179462 345470 179522 345478
rect 295609 345475 295675 345478
rect 179462 345410 180044 345470
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 296621 343498 296687 343501
rect 292836 343496 296687 343498
rect 292836 343440 296626 343496
rect 296682 343440 296687 343496
rect 292836 343438 296687 343440
rect 296621 343435 296687 343438
rect 179462 343370 180044 343430
rect 179462 343365 179522 343370
rect 179413 343360 179522 343365
rect 179413 343304 179418 343360
rect 179474 343304 179522 343360
rect 179413 343302 179522 343304
rect 179413 343299 179479 343302
rect 49509 341458 49575 341461
rect 125726 341458 125732 341460
rect 49509 341456 125732 341458
rect 49509 341400 49514 341456
rect 49570 341400 125732 341456
rect 49509 341398 125732 341400
rect 49509 341395 49575 341398
rect 125726 341396 125732 341398
rect 125796 341458 125802 341460
rect 126881 341458 126947 341461
rect 125796 341456 126947 341458
rect 125796 341400 126886 341456
rect 126942 341400 126947 341456
rect 125796 341398 126947 341400
rect 125796 341396 125802 341398
rect 126881 341395 126947 341398
rect 179505 341390 179571 341393
rect 179505 341388 180044 341390
rect 179505 341332 179510 341388
rect 179566 341332 180044 341388
rect 179505 341330 180044 341332
rect 179505 341327 179571 341330
rect 295609 340778 295675 340781
rect 292836 340776 295675 340778
rect 292836 340720 295614 340776
rect 295670 340720 295675 340776
rect 292836 340718 295675 340720
rect 295609 340715 295675 340718
rect 179462 339290 180044 339350
rect 176326 339220 176332 339284
rect 176396 339282 176402 339284
rect 179462 339282 179522 339290
rect 176396 339222 179522 339282
rect 176396 339220 176402 339222
rect 295609 338738 295675 338741
rect 292836 338736 295675 338738
rect 292836 338680 295614 338736
rect 295670 338680 295675 338736
rect 292836 338678 295675 338680
rect 295609 338675 295675 338678
rect 583520 338452 584960 338692
rect 294137 336698 294203 336701
rect 292836 336696 294203 336698
rect 292836 336640 294142 336696
rect 294198 336640 294203 336696
rect 292836 336638 294203 336640
rect 294137 336635 294203 336638
rect 179462 336570 180044 336630
rect 176561 336562 176627 336565
rect 179462 336562 179522 336570
rect 176561 336560 179522 336562
rect 176561 336504 176566 336560
rect 176622 336504 179522 336560
rect 176561 336502 179522 336504
rect 176561 336499 176627 336502
rect 293217 334658 293283 334661
rect 292836 334656 293283 334658
rect 292836 334600 293222 334656
rect 293278 334600 293283 334656
rect 292836 334598 293283 334600
rect 293217 334595 293283 334598
rect 179462 334530 180044 334590
rect 176653 334522 176719 334525
rect 179462 334522 179522 334530
rect 176653 334520 179522 334522
rect 176653 334464 176658 334520
rect 176714 334464 179522 334520
rect 176653 334462 179522 334464
rect 176653 334459 176719 334462
rect 176469 332618 176535 332621
rect 176469 332616 179890 332618
rect 176469 332560 176474 332616
rect 176530 332560 179890 332616
rect 176469 332558 179890 332560
rect 176469 332555 176535 332558
rect 179830 332550 179890 332558
rect 179830 332490 180044 332550
rect -960 332196 480 332436
rect 294045 331938 294111 331941
rect 292836 331936 294111 331938
rect 292836 331880 294050 331936
rect 294106 331880 294111 331936
rect 292836 331878 294111 331880
rect 294045 331875 294111 331878
rect 179462 330450 180044 330510
rect 176653 330442 176719 330445
rect 179462 330442 179522 330450
rect 176653 330440 179522 330442
rect 176653 330384 176658 330440
rect 176714 330384 179522 330440
rect 176653 330382 179522 330384
rect 176653 330379 176719 330382
rect 296897 329898 296963 329901
rect 292836 329896 296963 329898
rect 292836 329840 296902 329896
rect 296958 329840 296963 329896
rect 292836 329838 296963 329840
rect 296897 329835 296963 329838
rect 295517 327858 295583 327861
rect 292836 327856 295583 327858
rect 292836 327800 295522 327856
rect 295578 327800 295583 327856
rect 292836 327798 295583 327800
rect 295517 327795 295583 327798
rect 179462 327730 180044 327790
rect 59118 327660 59124 327724
rect 59188 327722 59194 327724
rect 139485 327722 139551 327725
rect 59188 327720 139551 327722
rect 59188 327664 139490 327720
rect 139546 327664 139551 327720
rect 59188 327662 139551 327664
rect 59188 327660 59194 327662
rect 139485 327659 139551 327662
rect 179270 327660 179276 327724
rect 179340 327722 179346 327724
rect 179462 327722 179522 327730
rect 179340 327662 179522 327722
rect 179340 327660 179346 327662
rect 176653 325818 176719 325821
rect 294045 325818 294111 325821
rect 176653 325816 179522 325818
rect 176653 325760 176658 325816
rect 176714 325760 179522 325816
rect 176653 325758 179522 325760
rect 292836 325816 294111 325818
rect 292836 325760 294050 325816
rect 294106 325760 294111 325816
rect 292836 325758 294111 325760
rect 176653 325755 176719 325758
rect 179462 325750 179522 325758
rect 294045 325755 294111 325758
rect 179462 325690 180044 325750
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 179462 323650 180044 323710
rect 176469 323642 176535 323645
rect 179462 323642 179522 323650
rect 176469 323640 179522 323642
rect 176469 323584 176474 323640
rect 176530 323584 179522 323640
rect 176469 323582 179522 323584
rect 176469 323579 176535 323582
rect 296621 323098 296687 323101
rect 292836 323096 296687 323098
rect 292836 323040 296626 323096
rect 296682 323040 296687 323096
rect 292836 323038 296687 323040
rect 296621 323035 296687 323038
rect 179462 321610 180044 321670
rect 175038 321540 175044 321604
rect 175108 321602 175114 321604
rect 179462 321602 179522 321610
rect 175108 321542 179522 321602
rect 175108 321540 175114 321542
rect 295425 321058 295491 321061
rect 292836 321056 295491 321058
rect 292836 321000 295430 321056
rect 295486 321000 295491 321056
rect 292836 320998 295491 321000
rect 295425 320995 295491 320998
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 295425 319018 295491 319021
rect 292836 319016 295491 319018
rect 292836 318960 295430 319016
rect 295486 318960 295491 319016
rect 292836 318958 295491 318960
rect 295425 318955 295491 318958
rect 179462 318890 180044 318950
rect 177665 318882 177731 318885
rect 179462 318882 179522 318890
rect 177665 318880 179522 318882
rect 177665 318824 177670 318880
rect 177726 318824 179522 318880
rect 177665 318822 179522 318824
rect 177665 318819 177731 318822
rect 295425 316978 295491 316981
rect 292836 316976 295491 316978
rect 292836 316920 295430 316976
rect 295486 316920 295491 316976
rect 292836 316918 295491 316920
rect 295425 316915 295491 316918
rect 179462 316850 180044 316910
rect 177573 316842 177639 316845
rect 179462 316842 179522 316850
rect 177573 316840 179522 316842
rect 177573 316784 177578 316840
rect 177634 316784 179522 316840
rect 177573 316782 179522 316784
rect 177573 316779 177639 316782
rect 176653 314938 176719 314941
rect 176653 314936 179522 314938
rect 176653 314880 176658 314936
rect 176714 314880 179522 314936
rect 176653 314878 179522 314880
rect 176653 314875 176719 314878
rect 179462 314870 179522 314878
rect 179462 314810 180044 314870
rect 49550 314740 49556 314804
rect 49620 314802 49626 314804
rect 59169 314802 59235 314805
rect 161974 314802 161980 314804
rect 49620 314800 161980 314802
rect 49620 314744 59174 314800
rect 59230 314744 161980 314800
rect 49620 314742 161980 314744
rect 49620 314740 49626 314742
rect 59169 314739 59235 314742
rect 161974 314740 161980 314742
rect 162044 314802 162050 314804
rect 162761 314802 162827 314805
rect 162044 314800 162827 314802
rect 162044 314744 162766 314800
rect 162822 314744 162827 314800
rect 162044 314742 162827 314744
rect 162044 314740 162050 314742
rect 162761 314739 162827 314742
rect 293125 314258 293191 314261
rect 293861 314258 293927 314261
rect 292836 314256 293927 314258
rect 292836 314200 293130 314256
rect 293186 314200 293866 314256
rect 293922 314200 293927 314256
rect 292836 314198 293927 314200
rect 293125 314195 293191 314198
rect 293861 314195 293927 314198
rect 176653 312898 176719 312901
rect 176653 312896 179522 312898
rect 176653 312840 176658 312896
rect 176714 312840 179522 312896
rect 176653 312838 179522 312840
rect 176653 312835 176719 312838
rect 179462 312830 179522 312838
rect 179462 312770 180044 312830
rect 294137 312218 294203 312221
rect 295374 312218 295380 312220
rect 292836 312216 295380 312218
rect 292836 312160 294142 312216
rect 294198 312160 295380 312216
rect 292836 312158 295380 312160
rect 294137 312155 294203 312158
rect 295374 312156 295380 312158
rect 295444 312156 295450 312220
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 295333 310178 295399 310181
rect 292836 310176 295399 310178
rect 292836 310120 295338 310176
rect 295394 310120 295399 310176
rect 292836 310118 295399 310120
rect 295333 310115 295399 310118
rect 179830 310050 180044 310110
rect 176653 310042 176719 310045
rect 177941 310042 178007 310045
rect 179830 310042 179890 310050
rect 176653 310040 179890 310042
rect 176653 309984 176658 310040
rect 176714 309984 177946 310040
rect 178002 309984 179890 310040
rect 176653 309982 179890 309984
rect 176653 309979 176719 309982
rect 177941 309979 178007 309982
rect 293166 309028 293172 309092
rect 293236 309090 293242 309092
rect 294229 309090 294295 309093
rect 293236 309088 294295 309090
rect 293236 309032 294234 309088
rect 294290 309032 294295 309088
rect 293236 309030 294295 309032
rect 293236 309028 293242 309030
rect 294229 309027 294295 309030
rect 295517 308138 295583 308141
rect 292836 308136 295583 308138
rect 292836 308080 295522 308136
rect 295578 308080 295583 308136
rect 292836 308078 295583 308080
rect 295517 308075 295583 308078
rect 179462 308010 180044 308070
rect 177941 308002 178007 308005
rect 179462 308002 179522 308010
rect 177941 308000 179522 308002
rect 177941 307944 177946 308000
rect 178002 307944 179522 308000
rect 177941 307942 179522 307944
rect 177941 307939 178007 307942
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 179830 305970 180044 306030
rect 177849 305962 177915 305965
rect 179830 305962 179890 305970
rect 177849 305960 179890 305962
rect 177849 305904 177854 305960
rect 177910 305904 179890 305960
rect 177849 305902 179890 305904
rect 177849 305899 177915 305902
rect 293902 305418 293908 305420
rect 292836 305358 293908 305418
rect 293902 305356 293908 305358
rect 293972 305356 293978 305420
rect 89713 305010 89779 305013
rect 90357 305010 90423 305013
rect 128854 305010 128860 305012
rect 89713 305008 128860 305010
rect 89713 304952 89718 305008
rect 89774 304952 90362 305008
rect 90418 304952 128860 305008
rect 89713 304950 128860 304952
rect 89713 304947 89779 304950
rect 90357 304947 90423 304950
rect 128854 304948 128860 304950
rect 128924 304948 128930 305012
rect 179462 303930 180044 303990
rect 176653 303922 176719 303925
rect 179462 303922 179522 303930
rect 176653 303920 179522 303922
rect 176653 303864 176658 303920
rect 176714 303864 179522 303920
rect 176653 303862 179522 303864
rect 176653 303859 176719 303862
rect 88977 303650 89043 303653
rect 148174 303650 148180 303652
rect 88977 303648 148180 303650
rect 88977 303592 88982 303648
rect 89038 303592 148180 303648
rect 88977 303590 148180 303592
rect 88977 303587 89043 303590
rect 148174 303588 148180 303590
rect 148244 303588 148250 303652
rect 292614 303452 292620 303516
rect 292684 303452 292690 303516
rect 292622 303348 292682 303452
rect 37181 301474 37247 301477
rect 124254 301474 124260 301476
rect 37181 301472 124260 301474
rect 37181 301416 37186 301472
rect 37242 301416 124260 301472
rect 37181 301414 124260 301416
rect 37181 301411 37247 301414
rect 124254 301412 124260 301414
rect 124324 301412 124330 301476
rect 143625 301474 143691 301477
rect 144678 301474 144684 301476
rect 143625 301472 144684 301474
rect 143625 301416 143630 301472
rect 143686 301416 144684 301472
rect 143625 301414 144684 301416
rect 143625 301411 143691 301414
rect 144678 301412 144684 301414
rect 144748 301412 144754 301476
rect 295333 301338 295399 301341
rect 292836 301336 295399 301338
rect 292836 301280 295338 301336
rect 295394 301280 295399 301336
rect 292836 301278 295399 301280
rect 295333 301275 295399 301278
rect 179462 301210 180044 301270
rect 73705 301202 73771 301205
rect 152406 301202 152412 301204
rect 73705 301200 152412 301202
rect 73705 301144 73710 301200
rect 73766 301144 152412 301200
rect 73705 301142 152412 301144
rect 73705 301139 73771 301142
rect 152406 301140 152412 301142
rect 152476 301140 152482 301204
rect 177849 301202 177915 301205
rect 179462 301202 179522 301210
rect 177849 301200 179522 301202
rect 177849 301144 177854 301200
rect 177910 301144 179522 301200
rect 177849 301142 179522 301144
rect 177849 301139 177915 301142
rect 109125 301066 109191 301069
rect 110321 301066 110387 301069
rect 138606 301066 138612 301068
rect 109125 301064 138612 301066
rect 109125 301008 109130 301064
rect 109186 301008 110326 301064
rect 110382 301008 138612 301064
rect 109125 301006 138612 301008
rect 109125 301003 109191 301006
rect 110321 301003 110387 301006
rect 138606 301004 138612 301006
rect 138676 301004 138682 301068
rect 107653 300794 107719 300797
rect 108941 300794 109007 300797
rect 107653 300792 109007 300794
rect 107653 300736 107658 300792
rect 107714 300736 108946 300792
rect 109002 300736 109007 300792
rect 107653 300734 109007 300736
rect 107653 300731 107719 300734
rect 108941 300731 109007 300734
rect 108941 299570 109007 299573
rect 130326 299570 130332 299572
rect 108941 299568 130332 299570
rect 108941 299512 108946 299568
rect 109002 299512 130332 299568
rect 108941 299510 130332 299512
rect 108941 299507 109007 299510
rect 130326 299508 130332 299510
rect 130396 299508 130402 299572
rect 176653 299298 176719 299301
rect 295333 299298 295399 299301
rect 176653 299296 179522 299298
rect 176653 299240 176658 299296
rect 176714 299240 179522 299296
rect 176653 299238 179522 299240
rect 292836 299296 295399 299298
rect 292836 299240 295338 299296
rect 295394 299240 295399 299296
rect 292836 299238 295399 299240
rect 176653 299235 176719 299238
rect 179462 299230 179522 299238
rect 295333 299235 295399 299238
rect 179462 299170 180044 299230
rect 112437 298890 112503 298893
rect 118969 298890 119035 298893
rect 112437 298888 119035 298890
rect 112437 298832 112442 298888
rect 112498 298832 118974 298888
rect 119030 298832 119035 298888
rect 112437 298830 119035 298832
rect 112437 298827 112503 298830
rect 118969 298827 119035 298830
rect 69054 298692 69060 298756
rect 69124 298754 69130 298756
rect 149053 298754 149119 298757
rect 162209 298754 162275 298757
rect 69124 298752 162275 298754
rect 69124 298696 149058 298752
rect 149114 298696 162214 298752
rect 162270 298696 162275 298752
rect 69124 298694 162275 298696
rect 69124 298692 69130 298694
rect 149053 298691 149119 298694
rect 162209 298691 162275 298694
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 176653 297258 176719 297261
rect 176653 297256 179522 297258
rect 176653 297200 176658 297256
rect 176714 297200 179522 297256
rect 176653 297198 179522 297200
rect 176653 297195 176719 297198
rect 179462 297190 179522 297198
rect 179462 297130 180044 297190
rect 103421 296986 103487 296989
rect 104341 296986 104407 296989
rect 153694 296986 153700 296988
rect 103421 296984 153700 296986
rect 103421 296928 103426 296984
rect 103482 296928 104346 296984
rect 104402 296928 153700 296984
rect 103421 296926 153700 296928
rect 103421 296923 103487 296926
rect 104341 296923 104407 296926
rect 153694 296924 153700 296926
rect 153764 296924 153770 296988
rect 67541 296850 67607 296853
rect 157977 296850 158043 296853
rect 67541 296848 158043 296850
rect 67541 296792 67546 296848
rect 67602 296792 157982 296848
rect 158038 296792 158043 296848
rect 67541 296790 158043 296792
rect 67541 296787 67607 296790
rect 157977 296787 158043 296790
rect 295517 296578 295583 296581
rect 292836 296576 295583 296578
rect 292836 296520 295522 296576
rect 295578 296520 295583 296576
rect 292836 296518 295583 296520
rect 295517 296515 295583 296518
rect 117681 295626 117747 295629
rect 118601 295626 118667 295629
rect 169702 295626 169708 295628
rect 117681 295624 169708 295626
rect 117681 295568 117686 295624
rect 117742 295568 118606 295624
rect 118662 295568 169708 295624
rect 117681 295566 169708 295568
rect 117681 295563 117747 295566
rect 118601 295563 118667 295566
rect 169702 295564 169708 295566
rect 169772 295564 169778 295628
rect 103513 295490 103579 295493
rect 104157 295490 104223 295493
rect 160686 295490 160692 295492
rect 103513 295488 160692 295490
rect 103513 295432 103518 295488
rect 103574 295432 104162 295488
rect 104218 295432 160692 295488
rect 103513 295430 160692 295432
rect 103513 295427 103579 295430
rect 104157 295427 104223 295430
rect 160686 295428 160692 295430
rect 160756 295428 160762 295492
rect 71773 295354 71839 295357
rect 171869 295354 171935 295357
rect 172421 295354 172487 295357
rect 71773 295352 172487 295354
rect 71773 295296 71778 295352
rect 71834 295296 171874 295352
rect 171930 295296 172426 295352
rect 172482 295296 172487 295352
rect 71773 295294 172487 295296
rect 71773 295291 71839 295294
rect 73846 295221 73906 295294
rect 171869 295291 171935 295294
rect 172421 295291 172487 295294
rect 73846 295216 73955 295221
rect 73846 295160 73894 295216
rect 73950 295160 73955 295216
rect 73846 295158 73955 295160
rect 73889 295155 73955 295158
rect 176653 295218 176719 295221
rect 176653 295216 179522 295218
rect 176653 295160 176658 295216
rect 176714 295160 179522 295216
rect 176653 295158 179522 295160
rect 176653 295155 176719 295158
rect 179462 295150 179522 295158
rect 179462 295090 180044 295150
rect 64689 294540 64755 294541
rect 64638 294476 64644 294540
rect 64708 294538 64755 294540
rect 75821 294538 75887 294541
rect 76005 294538 76071 294541
rect 173566 294538 173572 294540
rect 64708 294536 64800 294538
rect 64750 294480 64800 294536
rect 64708 294478 64800 294480
rect 75821 294536 173572 294538
rect 75821 294480 75826 294536
rect 75882 294480 76010 294536
rect 76066 294480 173572 294536
rect 75821 294478 173572 294480
rect 64708 294476 64755 294478
rect 64689 294475 64755 294476
rect 75821 294475 75887 294478
rect 76005 294475 76071 294478
rect 173566 294476 173572 294478
rect 173636 294476 173642 294540
rect 295333 294538 295399 294541
rect 292836 294536 295399 294538
rect 292836 294480 295338 294536
rect 295394 294480 295399 294536
rect 292836 294478 295399 294480
rect 295333 294475 295399 294478
rect 78397 294266 78463 294269
rect 167821 294266 167887 294269
rect 78397 294264 167887 294266
rect 78397 294208 78402 294264
rect 78458 294208 167826 294264
rect 167882 294208 167887 294264
rect 78397 294206 167887 294208
rect 78397 294203 78463 294206
rect 167821 294203 167887 294206
rect 111885 294130 111951 294133
rect 141509 294130 141575 294133
rect 111885 294128 141575 294130
rect 111885 294072 111890 294128
rect 111946 294072 141514 294128
rect 141570 294072 141575 294128
rect 111885 294070 141575 294072
rect 111885 294067 111951 294070
rect 141509 294067 141575 294070
rect 173709 293994 173775 293997
rect 174486 293994 174492 293996
rect 173709 293992 174492 293994
rect 173709 293936 173714 293992
rect 173770 293936 174492 293992
rect 173709 293934 174492 293936
rect 173709 293931 173775 293934
rect 174486 293932 174492 293934
rect 174556 293932 174562 293996
rect -960 293178 480 293268
rect 2865 293178 2931 293181
rect -960 293176 2931 293178
rect -960 293120 2870 293176
rect 2926 293120 2931 293176
rect -960 293118 2931 293120
rect -960 293028 480 293118
rect 2865 293115 2931 293118
rect 68737 292906 68803 292909
rect 169109 292906 169175 292909
rect 68737 292904 169175 292906
rect 68737 292848 68742 292904
rect 68798 292848 169114 292904
rect 169170 292848 169175 292904
rect 68737 292846 169175 292848
rect 68737 292843 68803 292846
rect 169109 292843 169175 292846
rect 105537 292770 105603 292773
rect 106089 292770 106155 292773
rect 169293 292770 169359 292773
rect 105537 292768 169359 292770
rect 105537 292712 105542 292768
rect 105598 292712 106094 292768
rect 106150 292712 169298 292768
rect 169354 292712 169359 292768
rect 105537 292710 169359 292712
rect 105537 292707 105603 292710
rect 106089 292707 106155 292710
rect 169293 292707 169359 292710
rect 113817 292634 113883 292637
rect 122046 292634 122052 292636
rect 113817 292632 122052 292634
rect 113817 292576 113822 292632
rect 113878 292576 122052 292632
rect 113817 292574 122052 292576
rect 113817 292571 113883 292574
rect 122046 292572 122052 292574
rect 122116 292572 122122 292636
rect 295609 292498 295675 292501
rect 292836 292496 295675 292498
rect 292836 292440 295614 292496
rect 295670 292440 295675 292496
rect 292836 292438 295675 292440
rect 295609 292435 295675 292438
rect 179462 292370 180044 292430
rect 70485 292362 70551 292365
rect 179229 292362 179295 292365
rect 179462 292362 179522 292370
rect 70485 292360 70594 292362
rect 70485 292304 70490 292360
rect 70546 292304 70594 292360
rect 70485 292299 70594 292304
rect 179229 292360 179522 292362
rect 179229 292304 179234 292360
rect 179290 292304 179522 292360
rect 179229 292302 179522 292304
rect 179229 292299 179295 292302
rect 70534 291788 70594 292299
rect 117957 292090 118023 292093
rect 117957 292088 122850 292090
rect 117957 292032 117962 292088
rect 118018 292032 122850 292088
rect 117957 292030 122850 292032
rect 117957 292027 118023 292030
rect 119061 291954 119127 291957
rect 120022 291954 120028 291956
rect 119061 291952 120028 291954
rect 119061 291896 119066 291952
rect 119122 291896 120028 291952
rect 119061 291894 120028 291896
rect 119061 291891 119127 291894
rect 120022 291892 120028 291894
rect 120092 291892 120098 291956
rect 122790 291954 122850 292030
rect 142797 291954 142863 291957
rect 122790 291952 142863 291954
rect 122790 291896 142802 291952
rect 142858 291896 142863 291952
rect 122790 291894 142863 291896
rect 142797 291891 142863 291894
rect 121453 291818 121519 291821
rect 119876 291816 121519 291818
rect 119876 291760 121458 291816
rect 121514 291760 121519 291816
rect 119876 291758 121519 291760
rect 121453 291755 121519 291758
rect 67725 291138 67791 291141
rect 121637 291138 121703 291141
rect 67725 291136 70196 291138
rect 67725 291080 67730 291136
rect 67786 291080 70196 291136
rect 67725 291078 70196 291080
rect 119876 291136 121703 291138
rect 119876 291080 121642 291136
rect 121698 291080 121703 291136
rect 119876 291078 121703 291080
rect 67725 291075 67791 291078
rect 121637 291075 121703 291078
rect 67633 290458 67699 290461
rect 121453 290458 121519 290461
rect 67633 290456 70196 290458
rect 67633 290400 67638 290456
rect 67694 290400 70196 290456
rect 67633 290398 70196 290400
rect 119876 290456 121519 290458
rect 119876 290400 121458 290456
rect 121514 290400 121519 290456
rect 119876 290398 121519 290400
rect 67633 290395 67699 290398
rect 121453 290395 121519 290398
rect 124070 290396 124076 290460
rect 124140 290458 124146 290460
rect 166993 290458 167059 290461
rect 124140 290456 167059 290458
rect 124140 290400 166998 290456
rect 167054 290400 167059 290456
rect 124140 290398 167059 290400
rect 124140 290396 124146 290398
rect 166993 290395 167059 290398
rect 176653 290458 176719 290461
rect 295517 290458 295583 290461
rect 176653 290456 179522 290458
rect 176653 290400 176658 290456
rect 176714 290400 179522 290456
rect 176653 290398 179522 290400
rect 292836 290456 295583 290458
rect 292836 290400 295522 290456
rect 295578 290400 295583 290456
rect 292836 290398 295583 290400
rect 176653 290395 176719 290398
rect 179462 290390 179522 290398
rect 295517 290395 295583 290398
rect 179462 290330 180044 290390
rect 67725 289778 67791 289781
rect 67725 289776 70196 289778
rect 67725 289720 67730 289776
rect 67786 289720 70196 289776
rect 67725 289718 70196 289720
rect 67725 289715 67791 289718
rect 119846 289234 119906 289748
rect 129038 289234 129044 289236
rect 119846 289174 129044 289234
rect 129038 289172 129044 289174
rect 129108 289172 129114 289236
rect 67633 289098 67699 289101
rect 121453 289098 121519 289101
rect 67633 289096 70196 289098
rect 67633 289040 67638 289096
rect 67694 289040 70196 289096
rect 67633 289038 70196 289040
rect 119876 289096 121519 289098
rect 119876 289040 121458 289096
rect 121514 289040 121519 289096
rect 119876 289038 121519 289040
rect 67633 289035 67699 289038
rect 121453 289035 121519 289038
rect 121637 288418 121703 288421
rect 119876 288416 121703 288418
rect 70534 288148 70594 288388
rect 119876 288360 121642 288416
rect 121698 288360 121703 288416
rect 119876 288358 121703 288360
rect 121637 288355 121703 288358
rect 176653 288418 176719 288421
rect 176653 288416 179522 288418
rect 176653 288360 176658 288416
rect 176714 288360 179522 288416
rect 176653 288358 179522 288360
rect 176653 288355 176719 288358
rect 179462 288350 179522 288358
rect 179462 288290 180044 288350
rect 70526 288084 70532 288148
rect 70596 288084 70602 288148
rect 67633 287738 67699 287741
rect 121453 287738 121519 287741
rect 293125 287738 293191 287741
rect 67633 287736 70196 287738
rect 67633 287680 67638 287736
rect 67694 287680 70196 287736
rect 67633 287678 70196 287680
rect 119876 287736 121519 287738
rect 119876 287680 121458 287736
rect 121514 287680 121519 287736
rect 119876 287678 121519 287680
rect 292836 287736 293191 287738
rect 292836 287680 293130 287736
rect 293186 287680 293191 287736
rect 292836 287678 293191 287680
rect 67633 287675 67699 287678
rect 121453 287675 121519 287678
rect 293125 287675 293191 287678
rect 67817 287058 67883 287061
rect 124254 287058 124260 287060
rect 67817 287056 70196 287058
rect 67817 287000 67822 287056
rect 67878 287000 70196 287056
rect 67817 286998 70196 287000
rect 119876 286998 124260 287058
rect 67817 286995 67883 286998
rect 124254 286996 124260 286998
rect 124324 286996 124330 287060
rect 124254 286588 124260 286652
rect 124324 286650 124330 286652
rect 124397 286650 124463 286653
rect 124324 286648 124463 286650
rect 124324 286592 124402 286648
rect 124458 286592 124463 286648
rect 124324 286590 124463 286592
rect 124324 286588 124330 286590
rect 124397 286587 124463 286590
rect 67725 286378 67791 286381
rect 120073 286378 120139 286381
rect 67725 286376 70196 286378
rect 67725 286320 67730 286376
rect 67786 286320 70196 286376
rect 67725 286318 70196 286320
rect 119876 286376 120139 286378
rect 119876 286320 120078 286376
rect 120134 286320 120139 286376
rect 119876 286318 120139 286320
rect 67725 286315 67791 286318
rect 120073 286315 120139 286318
rect 179462 286250 180044 286310
rect 179321 286242 179387 286245
rect 179462 286242 179522 286250
rect 161430 286240 179522 286242
rect 161430 286184 179326 286240
rect 179382 286184 179522 286240
rect 161430 286182 179522 286184
rect 120574 285908 120580 285972
rect 120644 285970 120650 285972
rect 161430 285970 161490 286182
rect 179321 286179 179387 286182
rect 120644 285910 161490 285970
rect 120644 285908 120650 285910
rect 69105 285698 69171 285701
rect 125726 285698 125732 285700
rect 69105 285696 70196 285698
rect 69105 285640 69110 285696
rect 69166 285640 70196 285696
rect 69105 285638 70196 285640
rect 119876 285638 125732 285698
rect 69105 285635 69171 285638
rect 125726 285636 125732 285638
rect 125796 285636 125802 285700
rect 295425 285698 295491 285701
rect 292836 285696 295491 285698
rect 292836 285640 295430 285696
rect 295486 285640 295491 285696
rect 292836 285638 295491 285640
rect 295425 285635 295491 285638
rect 583520 285276 584960 285516
rect 68737 285018 68803 285021
rect 121453 285018 121519 285021
rect 68737 285016 70196 285018
rect 68737 284960 68742 285016
rect 68798 284960 70196 285016
rect 68737 284958 70196 284960
rect 119876 285016 121519 285018
rect 119876 284960 121458 285016
rect 121514 284960 121519 285016
rect 119876 284958 121519 284960
rect 68737 284955 68803 284958
rect 121453 284955 121519 284958
rect 39849 284338 39915 284341
rect 53833 284338 53899 284341
rect 54334 284338 54340 284340
rect 39849 284336 54340 284338
rect 39849 284280 39854 284336
rect 39910 284280 53838 284336
rect 53894 284280 54340 284336
rect 39849 284278 54340 284280
rect 39849 284275 39915 284278
rect 53833 284275 53899 284278
rect 54334 284276 54340 284278
rect 54404 284276 54410 284340
rect 67633 284338 67699 284341
rect 121545 284338 121611 284341
rect 67633 284336 70196 284338
rect 67633 284280 67638 284336
rect 67694 284280 70196 284336
rect 67633 284278 70196 284280
rect 119876 284336 121611 284338
rect 119876 284280 121550 284336
rect 121606 284280 121611 284336
rect 119876 284278 121611 284280
rect 67633 284275 67699 284278
rect 121545 284275 121611 284278
rect 67725 283658 67791 283661
rect 176653 283658 176719 283661
rect 295425 283658 295491 283661
rect 67725 283656 70196 283658
rect 67725 283600 67730 283656
rect 67786 283600 70196 283656
rect 176653 283656 179522 283658
rect 67725 283598 70196 283600
rect 67725 283595 67791 283598
rect 119654 283324 119660 283388
rect 119724 283324 119730 283388
rect 67633 282978 67699 282981
rect 119662 282978 119722 283324
rect 119846 283250 119906 283628
rect 176653 283600 176658 283656
rect 176714 283600 179522 283656
rect 176653 283598 179522 283600
rect 292836 283656 295491 283658
rect 292836 283600 295430 283656
rect 295486 283600 295491 283656
rect 292836 283598 295491 283600
rect 176653 283595 176719 283598
rect 179462 283590 179522 283598
rect 295425 283595 295491 283598
rect 179462 283530 180044 283590
rect 126094 283250 126100 283252
rect 119846 283190 126100 283250
rect 126094 283188 126100 283190
rect 126164 283188 126170 283252
rect 121453 282978 121519 282981
rect 67633 282976 70196 282978
rect 67633 282920 67638 282976
rect 67694 282920 70196 282976
rect 119662 282976 121519 282978
rect 119662 282948 121458 282976
rect 67633 282918 70196 282920
rect 119692 282920 121458 282948
rect 121514 282920 121519 282976
rect 119692 282918 121519 282920
rect 67633 282915 67699 282918
rect 121453 282915 121519 282918
rect 121545 282298 121611 282301
rect 119876 282296 121611 282298
rect 119876 282240 121550 282296
rect 121606 282240 121611 282296
rect 119876 282238 121611 282240
rect 121545 282235 121611 282238
rect 292614 281692 292620 281756
rect 292684 281754 292690 281756
rect 292684 281694 292866 281754
rect 292684 281692 292690 281694
rect 68645 281618 68711 281621
rect 121453 281618 121519 281621
rect 68645 281616 70196 281618
rect 68645 281560 68650 281616
rect 68706 281560 70196 281616
rect 68645 281558 70196 281560
rect 119876 281616 121519 281618
rect 119876 281560 121458 281616
rect 121514 281560 121519 281616
rect 119876 281558 121519 281560
rect 68645 281555 68711 281558
rect 121453 281555 121519 281558
rect 176653 281618 176719 281621
rect 292806 281618 292866 281694
rect 295425 281618 295491 281621
rect 176653 281616 179522 281618
rect 176653 281560 176658 281616
rect 176714 281560 179522 281616
rect 292806 281616 295491 281618
rect 292806 281588 295430 281616
rect 176653 281558 179522 281560
rect 292836 281560 295430 281588
rect 295486 281560 295491 281616
rect 292836 281558 295491 281560
rect 176653 281555 176719 281558
rect 179462 281550 179522 281558
rect 295425 281555 295491 281558
rect 179462 281490 180044 281550
rect 67633 280938 67699 280941
rect 120165 280938 120231 280941
rect 122097 280938 122163 280941
rect 67633 280936 70196 280938
rect 67633 280880 67638 280936
rect 67694 280880 70196 280936
rect 67633 280878 70196 280880
rect 119876 280936 122163 280938
rect 119876 280880 120170 280936
rect 120226 280880 122102 280936
rect 122158 280880 122163 280936
rect 119876 280878 122163 280880
rect 67633 280875 67699 280878
rect 120165 280875 120231 280878
rect 122097 280875 122163 280878
rect 67633 280258 67699 280261
rect 121453 280258 121519 280261
rect 67633 280256 70196 280258
rect -960 279972 480 280212
rect 67633 280200 67638 280256
rect 67694 280200 70196 280256
rect 67633 280198 70196 280200
rect 119876 280256 121519 280258
rect 119876 280200 121458 280256
rect 121514 280200 121519 280256
rect 119876 280198 121519 280200
rect 67633 280195 67699 280198
rect 121453 280195 121519 280198
rect 67633 279578 67699 279581
rect 122741 279578 122807 279581
rect 67633 279576 70196 279578
rect 67633 279520 67638 279576
rect 67694 279520 70196 279576
rect 67633 279518 70196 279520
rect 119876 279576 122807 279578
rect 119876 279520 122746 279576
rect 122802 279520 122807 279576
rect 119876 279518 122807 279520
rect 67633 279515 67699 279518
rect 122741 279515 122807 279518
rect 176745 279578 176811 279581
rect 179086 279578 179092 279580
rect 176745 279576 179092 279578
rect 176745 279520 176750 279576
rect 176806 279520 179092 279576
rect 176745 279518 179092 279520
rect 176745 279515 176811 279518
rect 179086 279516 179092 279518
rect 179156 279578 179162 279580
rect 179156 279518 179890 279578
rect 179156 279516 179162 279518
rect 179830 279510 179890 279518
rect 179830 279450 180044 279510
rect 67725 278898 67791 278901
rect 121453 278898 121519 278901
rect 295425 278898 295491 278901
rect 67725 278896 70196 278898
rect 67725 278840 67730 278896
rect 67786 278840 70196 278896
rect 67725 278838 70196 278840
rect 119876 278896 121519 278898
rect 119876 278840 121458 278896
rect 121514 278840 121519 278896
rect 119876 278838 121519 278840
rect 292836 278896 295491 278898
rect 292836 278840 295430 278896
rect 295486 278840 295491 278896
rect 292836 278838 295491 278840
rect 67725 278835 67791 278838
rect 121453 278835 121519 278838
rect 295425 278835 295491 278838
rect 121637 278762 121703 278765
rect 122281 278762 122347 278765
rect 120214 278760 122347 278762
rect 120214 278704 121642 278760
rect 121698 278704 122286 278760
rect 122342 278704 122347 278760
rect 120214 278702 122347 278704
rect 120214 278626 120274 278702
rect 121637 278699 121703 278702
rect 122281 278699 122347 278702
rect 119846 278566 120274 278626
rect 67633 278218 67699 278221
rect 67633 278216 70196 278218
rect 67633 278160 67638 278216
rect 67694 278160 70196 278216
rect 119846 278188 119906 278566
rect 67633 278158 70196 278160
rect 67633 278155 67699 278158
rect 67633 277538 67699 277541
rect 121545 277538 121611 277541
rect 67633 277536 70196 277538
rect 67633 277480 67638 277536
rect 67694 277480 70196 277536
rect 67633 277478 70196 277480
rect 119876 277536 121611 277538
rect 119876 277480 121550 277536
rect 121606 277480 121611 277536
rect 119876 277478 121611 277480
rect 67633 277475 67699 277478
rect 121545 277475 121611 277478
rect 176653 277538 176719 277541
rect 176653 277536 179522 277538
rect 176653 277480 176658 277536
rect 176714 277480 179522 277536
rect 176653 277478 179522 277480
rect 176653 277475 176719 277478
rect 179462 277470 179522 277478
rect 179462 277410 180044 277470
rect 67725 276858 67791 276861
rect 121453 276858 121519 276861
rect 295425 276858 295491 276861
rect 67725 276856 70196 276858
rect 67725 276800 67730 276856
rect 67786 276800 70196 276856
rect 67725 276798 70196 276800
rect 119876 276856 121519 276858
rect 119876 276800 121458 276856
rect 121514 276800 121519 276856
rect 119876 276798 121519 276800
rect 292836 276856 295491 276858
rect 292836 276800 295430 276856
rect 295486 276800 295491 276856
rect 292836 276798 295491 276800
rect 67725 276795 67791 276798
rect 121453 276795 121519 276798
rect 295425 276795 295491 276798
rect 67633 276178 67699 276181
rect 67633 276176 70196 276178
rect 67633 276120 67638 276176
rect 67694 276120 70196 276176
rect 67633 276118 70196 276120
rect 119876 276118 122850 276178
rect 67633 276115 67699 276118
rect 122790 276042 122850 276118
rect 166390 276042 166396 276044
rect 122790 275982 166396 276042
rect 166390 275980 166396 275982
rect 166460 275980 166466 276044
rect 68185 275498 68251 275501
rect 68921 275498 68987 275501
rect 121453 275498 121519 275501
rect 68185 275496 70196 275498
rect 68185 275440 68190 275496
rect 68246 275440 68926 275496
rect 68982 275440 70196 275496
rect 68185 275438 70196 275440
rect 119876 275496 121519 275498
rect 119876 275440 121458 275496
rect 121514 275440 121519 275496
rect 119876 275438 121519 275440
rect 68185 275435 68251 275438
rect 68921 275435 68987 275438
rect 121453 275435 121519 275438
rect 67633 274818 67699 274821
rect 121545 274818 121611 274821
rect 67633 274816 70196 274818
rect 67633 274760 67638 274816
rect 67694 274760 70196 274816
rect 67633 274758 70196 274760
rect 119876 274816 121611 274818
rect 119876 274760 121550 274816
rect 121606 274760 121611 274816
rect 119876 274758 121611 274760
rect 67633 274755 67699 274758
rect 121545 274755 121611 274758
rect 176653 274818 176719 274821
rect 295425 274818 295491 274821
rect 176653 274816 179522 274818
rect 176653 274760 176658 274816
rect 176714 274760 179522 274816
rect 176653 274758 179522 274760
rect 292836 274816 295491 274818
rect 292836 274760 295430 274816
rect 295486 274760 295491 274816
rect 292836 274758 295491 274760
rect 176653 274755 176719 274758
rect 179462 274750 179522 274758
rect 295425 274755 295491 274758
rect 179462 274690 180044 274750
rect 68001 274138 68067 274141
rect 69105 274138 69171 274141
rect 121453 274138 121519 274141
rect 68001 274136 70196 274138
rect 68001 274080 68006 274136
rect 68062 274080 69110 274136
rect 69166 274080 70196 274136
rect 68001 274078 70196 274080
rect 119876 274136 121519 274138
rect 119876 274080 121458 274136
rect 121514 274080 121519 274136
rect 119876 274078 121519 274080
rect 68001 274075 68067 274078
rect 69105 274075 69171 274078
rect 121453 274075 121519 274078
rect 67817 273458 67883 273461
rect 121453 273458 121519 273461
rect 67817 273456 70196 273458
rect 67817 273400 67822 273456
rect 67878 273400 70196 273456
rect 67817 273398 70196 273400
rect 119876 273456 121519 273458
rect 119876 273400 121458 273456
rect 121514 273400 121519 273456
rect 119876 273398 121519 273400
rect 67817 273395 67883 273398
rect 121453 273395 121519 273398
rect 67633 272778 67699 272781
rect 121453 272778 121519 272781
rect 295425 272778 295491 272781
rect 67633 272776 70196 272778
rect 67633 272720 67638 272776
rect 67694 272720 70196 272776
rect 67633 272718 70196 272720
rect 119876 272776 121519 272778
rect 119876 272720 121458 272776
rect 121514 272720 121519 272776
rect 119876 272718 121519 272720
rect 292836 272776 295491 272778
rect 292836 272720 295430 272776
rect 295486 272720 295491 272776
rect 292836 272718 295491 272720
rect 67633 272715 67699 272718
rect 121453 272715 121519 272718
rect 295425 272715 295491 272718
rect 179462 272650 180044 272710
rect 145741 272642 145807 272645
rect 149646 272642 149652 272644
rect 145741 272640 149652 272642
rect 145741 272584 145746 272640
rect 145802 272584 149652 272640
rect 145741 272582 149652 272584
rect 145741 272579 145807 272582
rect 149646 272580 149652 272582
rect 149716 272580 149722 272644
rect 176653 272642 176719 272645
rect 179462 272642 179522 272650
rect 176653 272640 179522 272642
rect 176653 272584 176658 272640
rect 176714 272584 179522 272640
rect 176653 272582 179522 272584
rect 176653 272579 176719 272582
rect 582465 272234 582531 272237
rect 583520 272234 584960 272324
rect 582465 272232 584960 272234
rect 582465 272176 582470 272232
rect 582526 272176 584960 272232
rect 582465 272174 584960 272176
rect 582465 272171 582531 272174
rect 67817 272098 67883 272101
rect 122373 272098 122439 272101
rect 67817 272096 70196 272098
rect 67817 272040 67822 272096
rect 67878 272040 70196 272096
rect 67817 272038 70196 272040
rect 119876 272096 122439 272098
rect 119876 272040 122378 272096
rect 122434 272040 122439 272096
rect 583520 272084 584960 272174
rect 119876 272038 122439 272040
rect 67817 272035 67883 272038
rect 122373 272035 122439 272038
rect 54937 271826 55003 271829
rect 55622 271826 55628 271828
rect 54937 271824 55628 271826
rect 54937 271768 54942 271824
rect 54998 271768 55628 271824
rect 54937 271766 55628 271768
rect 54937 271763 55003 271766
rect 55622 271764 55628 271766
rect 55692 271764 55698 271828
rect 67725 271418 67791 271421
rect 121453 271418 121519 271421
rect 67725 271416 70196 271418
rect 67725 271360 67730 271416
rect 67786 271360 70196 271416
rect 67725 271358 70196 271360
rect 119876 271416 121519 271418
rect 119876 271360 121458 271416
rect 121514 271360 121519 271416
rect 119876 271358 121519 271360
rect 67725 271355 67791 271358
rect 121453 271355 121519 271358
rect 67633 270738 67699 270741
rect 67633 270736 70196 270738
rect 67633 270680 67638 270736
rect 67694 270680 70196 270736
rect 67633 270678 70196 270680
rect 67633 270675 67699 270678
rect 179462 270610 180044 270670
rect 177757 270602 177823 270605
rect 179462 270602 179522 270610
rect 177757 270600 179522 270602
rect 177757 270544 177762 270600
rect 177818 270544 179522 270600
rect 177757 270542 179522 270544
rect 177757 270539 177823 270542
rect 67725 270058 67791 270061
rect 121453 270058 121519 270061
rect 295425 270058 295491 270061
rect 67725 270056 70196 270058
rect 67725 270000 67730 270056
rect 67786 270000 70196 270056
rect 67725 269998 70196 270000
rect 119876 270056 121519 270058
rect 119876 270000 121458 270056
rect 121514 270000 121519 270056
rect 119876 269998 121519 270000
rect 292836 270056 295491 270058
rect 292836 270000 295430 270056
rect 295486 270000 295491 270056
rect 292836 269998 295491 270000
rect 67725 269995 67791 269998
rect 121453 269995 121519 269998
rect 295425 269995 295491 269998
rect 67633 269378 67699 269381
rect 121545 269378 121611 269381
rect 67633 269376 70196 269378
rect 67633 269320 67638 269376
rect 67694 269320 70196 269376
rect 67633 269318 70196 269320
rect 119876 269376 121611 269378
rect 119876 269320 121550 269376
rect 121606 269320 121611 269376
rect 119876 269318 121611 269320
rect 67633 269315 67699 269318
rect 121545 269315 121611 269318
rect 67725 268698 67791 268701
rect 121453 268698 121519 268701
rect 67725 268696 70196 268698
rect 67725 268640 67730 268696
rect 67786 268640 70196 268696
rect 67725 268638 70196 268640
rect 119876 268696 121519 268698
rect 119876 268640 121458 268696
rect 121514 268640 121519 268696
rect 119876 268638 121519 268640
rect 67725 268635 67791 268638
rect 121453 268635 121519 268638
rect 179462 268570 180044 268630
rect 179321 268562 179387 268565
rect 179462 268562 179522 268570
rect 179321 268560 179522 268562
rect 179321 268504 179326 268560
rect 179382 268504 179522 268560
rect 179321 268502 179522 268504
rect 179321 268499 179387 268502
rect 67633 268018 67699 268021
rect 121453 268018 121519 268021
rect 294229 268018 294295 268021
rect 67633 268016 70196 268018
rect 67633 267960 67638 268016
rect 67694 267960 70196 268016
rect 67633 267958 70196 267960
rect 119876 268016 121519 268018
rect 119876 267960 121458 268016
rect 121514 267960 121519 268016
rect 119876 267958 121519 267960
rect 292836 268016 294295 268018
rect 292836 267960 294234 268016
rect 294290 267960 294295 268016
rect 292836 267958 294295 267960
rect 67633 267955 67699 267958
rect 121453 267955 121519 267958
rect 294229 267955 294295 267958
rect 68645 267338 68711 267341
rect 121453 267338 121519 267341
rect 68645 267336 70196 267338
rect -960 267202 480 267292
rect 68645 267280 68650 267336
rect 68706 267280 70196 267336
rect 68645 267278 70196 267280
rect 119876 267336 121519 267338
rect 119876 267280 121458 267336
rect 121514 267280 121519 267336
rect 119876 267278 121519 267280
rect 68645 267275 68711 267278
rect 121453 267275 121519 267278
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 67541 266658 67607 266661
rect 121545 266658 121611 266661
rect 67541 266656 70196 266658
rect 67541 266600 67546 266656
rect 67602 266600 70196 266656
rect 67541 266598 70196 266600
rect 119876 266656 121611 266658
rect 119876 266600 121550 266656
rect 121606 266600 121611 266656
rect 119876 266598 121611 266600
rect 67541 266595 67607 266598
rect 121545 266595 121611 266598
rect 147581 266250 147647 266253
rect 122790 266248 147647 266250
rect 122790 266192 147586 266248
rect 147642 266192 147647 266248
rect 122790 266190 147647 266192
rect 68093 265978 68159 265981
rect 69197 265978 69263 265981
rect 122189 265978 122255 265981
rect 68093 265976 70196 265978
rect 68093 265920 68098 265976
rect 68154 265920 69202 265976
rect 69258 265920 70196 265976
rect 68093 265918 70196 265920
rect 119876 265976 122255 265978
rect 119876 265920 122194 265976
rect 122250 265920 122255 265976
rect 119876 265918 122255 265920
rect 68093 265915 68159 265918
rect 69197 265915 69263 265918
rect 122189 265915 122255 265918
rect 122790 265706 122850 266190
rect 147581 266187 147647 266190
rect 295425 265978 295491 265981
rect 292836 265976 295491 265978
rect 292836 265920 295430 265976
rect 295486 265920 295491 265976
rect 292836 265918 295491 265920
rect 295425 265915 295491 265918
rect 119846 265646 122850 265706
rect 179462 265850 180044 265910
rect 67633 265298 67699 265301
rect 67633 265296 70196 265298
rect 67633 265240 67638 265296
rect 67694 265240 70196 265296
rect 119846 265268 119906 265646
rect 147581 265570 147647 265573
rect 171726 265570 171732 265572
rect 147581 265568 171732 265570
rect 147581 265512 147586 265568
rect 147642 265512 171732 265568
rect 147581 265510 171732 265512
rect 147581 265507 147647 265510
rect 171726 265508 171732 265510
rect 171796 265508 171802 265572
rect 67633 265238 70196 265240
rect 67633 265235 67699 265238
rect 149646 264964 149652 265028
rect 149716 265026 149722 265028
rect 179462 265026 179522 265850
rect 149716 264966 179522 265026
rect 149716 264964 149722 264966
rect 67633 264618 67699 264621
rect 121453 264618 121519 264621
rect 67633 264616 70196 264618
rect 67633 264560 67638 264616
rect 67694 264560 70196 264616
rect 67633 264558 70196 264560
rect 119876 264616 121519 264618
rect 119876 264560 121458 264616
rect 121514 264560 121519 264616
rect 119876 264558 121519 264560
rect 67633 264555 67699 264558
rect 121453 264555 121519 264558
rect 68829 263938 68895 263941
rect 121545 263938 121611 263941
rect 295517 263938 295583 263941
rect 68829 263936 70196 263938
rect 68829 263880 68834 263936
rect 68890 263880 70196 263936
rect 68829 263878 70196 263880
rect 119876 263936 121611 263938
rect 119876 263880 121550 263936
rect 121606 263880 121611 263936
rect 119876 263878 121611 263880
rect 292836 263936 295583 263938
rect 292836 263880 295522 263936
rect 295578 263880 295583 263936
rect 292836 263878 295583 263880
rect 68829 263875 68895 263878
rect 121545 263875 121611 263878
rect 295517 263875 295583 263878
rect 179462 263810 180044 263870
rect 179137 263802 179203 263805
rect 179462 263802 179522 263810
rect 179137 263800 179522 263802
rect 179137 263744 179142 263800
rect 179198 263744 179522 263800
rect 179137 263742 179522 263744
rect 179137 263739 179203 263742
rect 67725 263258 67791 263261
rect 121453 263258 121519 263261
rect 67725 263256 70196 263258
rect 67725 263200 67730 263256
rect 67786 263200 70196 263256
rect 67725 263198 70196 263200
rect 119876 263256 121519 263258
rect 119876 263200 121458 263256
rect 121514 263200 121519 263256
rect 119876 263198 121519 263200
rect 67725 263195 67791 263198
rect 121453 263195 121519 263198
rect 67633 262578 67699 262581
rect 121453 262578 121519 262581
rect 67633 262576 70196 262578
rect 67633 262520 67638 262576
rect 67694 262520 70196 262576
rect 67633 262518 70196 262520
rect 119876 262576 121519 262578
rect 119876 262520 121458 262576
rect 121514 262520 121519 262576
rect 119876 262518 121519 262520
rect 67633 262515 67699 262518
rect 121453 262515 121519 262518
rect 177062 262108 177068 262172
rect 177132 262170 177138 262172
rect 179505 262170 179571 262173
rect 177132 262168 179571 262170
rect 177132 262112 179510 262168
rect 179566 262112 179571 262168
rect 177132 262110 179571 262112
rect 177132 262108 177138 262110
rect 179505 262107 179571 262110
rect 67633 261898 67699 261901
rect 120993 261898 121059 261901
rect 67633 261896 70196 261898
rect 67633 261840 67638 261896
rect 67694 261840 70196 261896
rect 67633 261838 70196 261840
rect 119876 261896 121059 261898
rect 119876 261840 120998 261896
rect 121054 261840 121059 261896
rect 119876 261838 121059 261840
rect 67633 261835 67699 261838
rect 120993 261835 121059 261838
rect 176653 261898 176719 261901
rect 176653 261896 179522 261898
rect 176653 261840 176658 261896
rect 176714 261840 179522 261896
rect 176653 261838 179522 261840
rect 176653 261835 176719 261838
rect 179462 261830 179522 261838
rect 179462 261770 180044 261830
rect 67725 261218 67791 261221
rect 121453 261218 121519 261221
rect 295425 261218 295491 261221
rect 67725 261216 70196 261218
rect 67725 261160 67730 261216
rect 67786 261160 70196 261216
rect 67725 261158 70196 261160
rect 119876 261216 121519 261218
rect 119876 261160 121458 261216
rect 121514 261160 121519 261216
rect 119876 261158 121519 261160
rect 292836 261216 295491 261218
rect 292836 261160 295430 261216
rect 295486 261160 295491 261216
rect 292836 261158 295491 261160
rect 67725 261155 67791 261158
rect 121453 261155 121519 261158
rect 295425 261155 295491 261158
rect 67633 260538 67699 260541
rect 121453 260538 121519 260541
rect 67633 260536 70196 260538
rect 67633 260480 67638 260536
rect 67694 260480 70196 260536
rect 67633 260478 70196 260480
rect 119876 260536 121519 260538
rect 119876 260480 121458 260536
rect 121514 260480 121519 260536
rect 119876 260478 121519 260480
rect 67633 260475 67699 260478
rect 121453 260475 121519 260478
rect 67725 259858 67791 259861
rect 121453 259858 121519 259861
rect 67725 259856 70196 259858
rect 67725 259800 67730 259856
rect 67786 259800 70196 259856
rect 67725 259798 70196 259800
rect 119876 259856 121519 259858
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 67725 259795 67791 259798
rect 121453 259795 121519 259798
rect 179462 259730 180044 259790
rect 177062 259660 177068 259724
rect 177132 259722 177138 259724
rect 179462 259722 179522 259730
rect 177132 259662 179522 259722
rect 177132 259660 177138 259662
rect 67725 259178 67791 259181
rect 122097 259178 122163 259181
rect 293217 259178 293283 259181
rect 67725 259176 70196 259178
rect 67725 259120 67730 259176
rect 67786 259120 70196 259176
rect 67725 259118 70196 259120
rect 119876 259176 122163 259178
rect 119876 259120 122102 259176
rect 122158 259120 122163 259176
rect 119876 259118 122163 259120
rect 292836 259176 293283 259178
rect 292836 259120 293222 259176
rect 293278 259120 293283 259176
rect 292836 259118 293283 259120
rect 67725 259115 67791 259118
rect 122097 259115 122163 259118
rect 293217 259115 293283 259118
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 67633 258498 67699 258501
rect 121453 258498 121519 258501
rect 67633 258496 70196 258498
rect 67633 258440 67638 258496
rect 67694 258440 70196 258496
rect 67633 258438 70196 258440
rect 119876 258496 121519 258498
rect 119876 258440 121458 258496
rect 121514 258440 121519 258496
rect 119876 258438 121519 258440
rect 67633 258435 67699 258438
rect 121453 258435 121519 258438
rect 67633 257818 67699 257821
rect 121545 257818 121611 257821
rect 67633 257816 70196 257818
rect 67633 257760 67638 257816
rect 67694 257760 70196 257816
rect 67633 257758 70196 257760
rect 119876 257816 121611 257818
rect 119876 257760 121550 257816
rect 121606 257760 121611 257816
rect 119876 257758 121611 257760
rect 67633 257755 67699 257758
rect 121545 257755 121611 257758
rect 121453 257138 121519 257141
rect 295374 257138 295380 257140
rect 119876 257136 121519 257138
rect 64454 256804 64460 256868
rect 64524 256866 64530 256868
rect 70166 256866 70226 257108
rect 119876 257080 121458 257136
rect 121514 257080 121519 257136
rect 119876 257078 121519 257080
rect 292836 257078 295380 257138
rect 121453 257075 121519 257078
rect 295374 257076 295380 257078
rect 295444 257076 295450 257140
rect 179462 257010 180044 257070
rect 176653 257002 176719 257005
rect 179462 257002 179522 257010
rect 176653 257000 179522 257002
rect 176653 256944 176658 257000
rect 176714 256944 179522 257000
rect 176653 256942 179522 256944
rect 176653 256939 176719 256942
rect 64524 256806 70226 256866
rect 64524 256804 64530 256806
rect 178769 256730 178835 256733
rect 179270 256730 179276 256732
rect 178769 256728 179276 256730
rect 178769 256672 178774 256728
rect 178830 256672 179276 256728
rect 178769 256670 179276 256672
rect 178769 256667 178835 256670
rect 179270 256668 179276 256670
rect 179340 256668 179346 256732
rect 67633 256458 67699 256461
rect 121545 256458 121611 256461
rect 67633 256456 70196 256458
rect 67633 256400 67638 256456
rect 67694 256400 70196 256456
rect 67633 256398 70196 256400
rect 119876 256456 121611 256458
rect 119876 256400 121550 256456
rect 121606 256400 121611 256456
rect 119876 256398 121611 256400
rect 67633 256395 67699 256398
rect 121545 256395 121611 256398
rect 122046 255852 122052 255916
rect 122116 255914 122122 255916
rect 149646 255914 149652 255916
rect 122116 255854 149652 255914
rect 122116 255852 122122 255854
rect 149646 255852 149652 255854
rect 149716 255852 149722 255916
rect 67909 255778 67975 255781
rect 68737 255778 68803 255781
rect 121453 255778 121519 255781
rect 67909 255776 70196 255778
rect 67909 255720 67914 255776
rect 67970 255720 68742 255776
rect 68798 255720 70196 255776
rect 67909 255718 70196 255720
rect 119876 255776 121519 255778
rect 119876 255720 121458 255776
rect 121514 255720 121519 255776
rect 119876 255718 121519 255720
rect 67909 255715 67975 255718
rect 68737 255715 68803 255718
rect 121453 255715 121519 255718
rect 172329 255236 172395 255237
rect 172278 255234 172284 255236
rect 172238 255174 172284 255234
rect 172348 255232 172395 255236
rect 172390 255176 172395 255232
rect 172278 255172 172284 255174
rect 172348 255172 172395 255176
rect 172329 255171 172395 255172
rect 67725 255098 67791 255101
rect 122373 255098 122439 255101
rect 295517 255098 295583 255101
rect 67725 255096 70196 255098
rect 67725 255040 67730 255096
rect 67786 255040 70196 255096
rect 67725 255038 70196 255040
rect 119876 255096 122439 255098
rect 119876 255040 122378 255096
rect 122434 255040 122439 255096
rect 119876 255038 122439 255040
rect 292836 255096 295583 255098
rect 292836 255040 295522 255096
rect 295578 255040 295583 255096
rect 292836 255038 295583 255040
rect 67725 255035 67791 255038
rect 122373 255035 122439 255038
rect 295517 255035 295583 255038
rect 179462 254970 180044 255030
rect 176653 254962 176719 254965
rect 179462 254962 179522 254970
rect 176653 254960 179522 254962
rect 176653 254904 176658 254960
rect 176714 254904 179522 254960
rect 176653 254902 179522 254904
rect 176653 254899 176719 254902
rect 67633 254418 67699 254421
rect 121453 254418 121519 254421
rect 67633 254416 70196 254418
rect 67633 254360 67638 254416
rect 67694 254360 70196 254416
rect 67633 254358 70196 254360
rect 119876 254416 121519 254418
rect 119876 254360 121458 254416
rect 121514 254360 121519 254416
rect 119876 254358 121519 254360
rect 67633 254355 67699 254358
rect 121453 254355 121519 254358
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 63125 254012 63191 254013
rect 63125 254008 63172 254012
rect 63236 254010 63242 254012
rect 63125 253952 63130 254008
rect 63125 253948 63172 253952
rect 63236 253950 63282 254010
rect 63236 253948 63242 253950
rect 63125 253947 63191 253948
rect 67633 253738 67699 253741
rect 121545 253738 121611 253741
rect 67633 253736 70196 253738
rect 67633 253680 67638 253736
rect 67694 253680 70196 253736
rect 67633 253678 70196 253680
rect 119876 253736 121611 253738
rect 119876 253680 121550 253736
rect 121606 253680 121611 253736
rect 119876 253678 121611 253680
rect 67633 253675 67699 253678
rect 121545 253675 121611 253678
rect 66846 252996 66852 253060
rect 66916 253058 66922 253060
rect 67398 253058 67404 253060
rect 66916 252998 67404 253058
rect 66916 252996 66922 252998
rect 67398 252996 67404 252998
rect 67468 253058 67474 253060
rect 121453 253058 121519 253061
rect 67468 252998 70196 253058
rect 119876 253056 121519 253058
rect 119876 253000 121458 253056
rect 121514 253000 121519 253056
rect 119876 252998 121519 253000
rect 67468 252996 67474 252998
rect 121453 252995 121519 252998
rect 179462 252930 180044 252990
rect 176653 252922 176719 252925
rect 179462 252922 179522 252930
rect 176653 252920 179522 252922
rect 176653 252864 176658 252920
rect 176714 252864 179522 252920
rect 176653 252862 179522 252864
rect 176653 252859 176719 252862
rect 63401 252516 63467 252517
rect 63350 252514 63356 252516
rect 63310 252454 63356 252514
rect 63420 252512 63467 252516
rect 63462 252456 63467 252512
rect 63350 252452 63356 252454
rect 63420 252452 63467 252456
rect 63401 252451 63467 252452
rect 69054 252316 69060 252380
rect 69124 252378 69130 252380
rect 121453 252378 121519 252381
rect 295517 252378 295583 252381
rect 69124 252318 70196 252378
rect 119876 252376 121519 252378
rect 119876 252320 121458 252376
rect 121514 252320 121519 252376
rect 119876 252318 121519 252320
rect 292836 252376 295583 252378
rect 292836 252320 295522 252376
rect 295578 252320 295583 252376
rect 292836 252318 295583 252320
rect 69124 252316 69130 252318
rect 121453 252315 121519 252318
rect 295517 252315 295583 252318
rect 67633 251698 67699 251701
rect 122189 251698 122255 251701
rect 67633 251696 70196 251698
rect 67633 251640 67638 251696
rect 67694 251640 70196 251696
rect 67633 251638 70196 251640
rect 119876 251696 122255 251698
rect 119876 251640 122194 251696
rect 122250 251640 122255 251696
rect 119876 251638 122255 251640
rect 67633 251635 67699 251638
rect 122189 251635 122255 251638
rect 67633 251018 67699 251021
rect 120165 251018 120231 251021
rect 120625 251018 120691 251021
rect 67633 251016 70196 251018
rect 67633 250960 67638 251016
rect 67694 250960 70196 251016
rect 67633 250958 70196 250960
rect 119876 251016 120691 251018
rect 119876 250960 120170 251016
rect 120226 250960 120630 251016
rect 120686 250960 120691 251016
rect 119876 250958 120691 250960
rect 67633 250955 67699 250958
rect 120165 250955 120231 250958
rect 120625 250955 120691 250958
rect 179462 250890 180044 250950
rect 176653 250882 176719 250885
rect 179462 250882 179522 250890
rect 176653 250880 179522 250882
rect 176653 250824 176658 250880
rect 176714 250824 179522 250880
rect 176653 250822 179522 250824
rect 176653 250819 176719 250822
rect 67541 250338 67607 250341
rect 121545 250338 121611 250341
rect 295517 250338 295583 250341
rect 67541 250336 70196 250338
rect 67541 250280 67546 250336
rect 67602 250280 70196 250336
rect 67541 250278 70196 250280
rect 119876 250336 121611 250338
rect 119876 250280 121550 250336
rect 121606 250280 121611 250336
rect 119876 250278 121611 250280
rect 292836 250336 295583 250338
rect 292836 250280 295522 250336
rect 295578 250280 295583 250336
rect 292836 250278 295583 250280
rect 67541 250275 67607 250278
rect 121545 250275 121611 250278
rect 295517 250275 295583 250278
rect 67633 249658 67699 249661
rect 121453 249658 121519 249661
rect 67633 249656 70196 249658
rect 67633 249600 67638 249656
rect 67694 249600 70196 249656
rect 67633 249598 70196 249600
rect 119876 249656 121519 249658
rect 119876 249600 121458 249656
rect 121514 249600 121519 249656
rect 119876 249598 121519 249600
rect 67633 249595 67699 249598
rect 121453 249595 121519 249598
rect 67633 248978 67699 248981
rect 122925 248978 122991 248981
rect 67633 248976 70196 248978
rect 67633 248920 67638 248976
rect 67694 248920 70196 248976
rect 67633 248918 70196 248920
rect 119876 248976 122991 248978
rect 119876 248920 122930 248976
rect 122986 248920 122991 248976
rect 119876 248918 122991 248920
rect 67633 248915 67699 248918
rect 122925 248915 122991 248918
rect 67725 248298 67791 248301
rect 121545 248298 121611 248301
rect 295006 248298 295012 248300
rect 67725 248296 70196 248298
rect 67725 248240 67730 248296
rect 67786 248240 70196 248296
rect 67725 248238 70196 248240
rect 119876 248296 121611 248298
rect 119876 248240 121550 248296
rect 121606 248240 121611 248296
rect 119876 248238 121611 248240
rect 292836 248238 295012 248298
rect 67725 248235 67791 248238
rect 121545 248235 121611 248238
rect 295006 248236 295012 248238
rect 295076 248236 295082 248300
rect 179462 248170 180044 248230
rect 179270 248100 179276 248164
rect 179340 248162 179346 248164
rect 179462 248162 179522 248170
rect 179340 248102 179522 248162
rect 179340 248100 179346 248102
rect 67633 247618 67699 247621
rect 121453 247618 121519 247621
rect 67633 247616 70196 247618
rect 67633 247560 67638 247616
rect 67694 247560 70196 247616
rect 67633 247558 70196 247560
rect 119876 247616 121519 247618
rect 119876 247560 121458 247616
rect 121514 247560 121519 247616
rect 119876 247558 121519 247560
rect 67633 247555 67699 247558
rect 121453 247555 121519 247558
rect 67633 246938 67699 246941
rect 121545 246938 121611 246941
rect 67633 246936 70196 246938
rect 67633 246880 67638 246936
rect 67694 246880 70196 246936
rect 67633 246878 70196 246880
rect 119876 246936 121611 246938
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 67633 246875 67699 246878
rect 121545 246875 121611 246878
rect 68185 246258 68251 246261
rect 121453 246258 121519 246261
rect 68185 246256 70196 246258
rect 68185 246200 68190 246256
rect 68246 246200 70196 246256
rect 68185 246198 70196 246200
rect 119876 246256 121519 246258
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 68185 246195 68251 246198
rect 121453 246195 121519 246198
rect 176653 246258 176719 246261
rect 295517 246260 295583 246261
rect 295517 246258 295564 246260
rect 176653 246256 179522 246258
rect 176653 246200 176658 246256
rect 176714 246200 179522 246256
rect 176653 246198 179522 246200
rect 292836 246256 295564 246258
rect 295628 246258 295634 246260
rect 292836 246200 295522 246256
rect 292836 246198 295564 246200
rect 176653 246195 176719 246198
rect 179462 246190 179522 246198
rect 295517 246196 295564 246198
rect 295628 246198 295710 246258
rect 295628 246196 295634 246198
rect 295517 246195 295583 246196
rect 179462 246130 180044 246190
rect 121453 245578 121519 245581
rect 119876 245576 121519 245578
rect 70166 245034 70226 245548
rect 119876 245520 121458 245576
rect 121514 245520 121519 245576
rect 119876 245518 121519 245520
rect 121453 245515 121519 245518
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 64830 244974 70226 245034
rect 61878 244428 61884 244492
rect 61948 244490 61954 244492
rect 64830 244490 64890 244974
rect 68185 244898 68251 244901
rect 121545 244898 121611 244901
rect 68185 244896 70196 244898
rect 68185 244840 68190 244896
rect 68246 244840 70196 244896
rect 68185 244838 70196 244840
rect 119876 244896 121611 244898
rect 119876 244840 121550 244896
rect 121606 244840 121611 244896
rect 119876 244838 121611 244840
rect 68185 244835 68251 244838
rect 121545 244835 121611 244838
rect 61948 244430 64890 244490
rect 61948 244428 61954 244430
rect 121453 244218 121519 244221
rect 119876 244216 121519 244218
rect 69657 243674 69723 243677
rect 70166 243674 70226 244188
rect 119876 244160 121458 244216
rect 121514 244160 121519 244216
rect 119876 244158 121519 244160
rect 121453 244155 121519 244158
rect 179597 244150 179663 244153
rect 179597 244148 180044 244150
rect 179597 244092 179602 244148
rect 179658 244092 180044 244148
rect 179597 244090 180044 244092
rect 179597 244087 179663 244090
rect 69657 243672 70226 243674
rect 69657 243616 69662 243672
rect 69718 243616 70226 243672
rect 69657 243614 70226 243616
rect 179413 243674 179479 243677
rect 179638 243674 179644 243676
rect 179413 243672 179644 243674
rect 179413 243616 179418 243672
rect 179474 243616 179644 243672
rect 179413 243614 179644 243616
rect 69657 243611 69723 243614
rect 179413 243611 179479 243614
rect 179638 243612 179644 243614
rect 179708 243612 179714 243676
rect 67633 243538 67699 243541
rect 67633 243536 70196 243538
rect 67633 243480 67638 243536
rect 67694 243480 70196 243536
rect 67633 243478 70196 243480
rect 67633 243475 67699 243478
rect 119846 242994 119906 243508
rect 144678 243476 144684 243540
rect 144748 243538 144754 243540
rect 166206 243538 166212 243540
rect 144748 243478 166212 243538
rect 144748 243476 144754 243478
rect 166206 243476 166212 243478
rect 166276 243476 166282 243540
rect 179505 243538 179571 243541
rect 179822 243538 179828 243540
rect 179505 243536 179828 243538
rect 179505 243480 179510 243536
rect 179566 243480 179828 243536
rect 179505 243478 179828 243480
rect 179505 243475 179571 243478
rect 179822 243476 179828 243478
rect 179892 243476 179898 243540
rect 296897 243538 296963 243541
rect 292836 243536 296963 243538
rect 292836 243480 296902 243536
rect 296958 243480 296963 243536
rect 292836 243478 296963 243480
rect 296897 243475 296963 243478
rect 146886 242994 146892 242996
rect 119846 242934 146892 242994
rect 146886 242932 146892 242934
rect 146956 242932 146962 242996
rect 67633 242858 67699 242861
rect 121453 242858 121519 242861
rect 67633 242856 70196 242858
rect 67633 242800 67638 242856
rect 67694 242800 70196 242856
rect 67633 242798 70196 242800
rect 119876 242856 121519 242858
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 67633 242795 67699 242798
rect 121453 242795 121519 242798
rect 67725 242178 67791 242181
rect 121545 242178 121611 242181
rect 67725 242176 70196 242178
rect 67725 242120 67730 242176
rect 67786 242120 70196 242176
rect 67725 242118 70196 242120
rect 119876 242176 121611 242178
rect 119876 242120 121550 242176
rect 121606 242120 121611 242176
rect 119876 242118 121611 242120
rect 67725 242115 67791 242118
rect 121545 242115 121611 242118
rect 179462 242050 180044 242110
rect 152406 241708 152412 241772
rect 152476 241770 152482 241772
rect 179462 241770 179522 242050
rect 152476 241710 179522 241770
rect 152476 241708 152482 241710
rect 67633 241498 67699 241501
rect 120073 241498 120139 241501
rect 67633 241496 70196 241498
rect 67633 241440 67638 241496
rect 67694 241440 70196 241496
rect 67633 241438 70196 241440
rect 119876 241496 120139 241498
rect 119876 241440 120078 241496
rect 120134 241440 120139 241496
rect 119876 241438 120139 241440
rect 67633 241435 67699 241438
rect 120073 241435 120139 241438
rect 126094 241436 126100 241500
rect 126164 241498 126170 241500
rect 165521 241498 165587 241501
rect 126164 241496 165587 241498
rect 126164 241440 165526 241496
rect 165582 241440 165587 241496
rect 126164 241438 165587 241440
rect 126164 241436 126170 241438
rect 165521 241435 165587 241438
rect 147121 241226 147187 241229
rect 292806 241226 292866 241468
rect 293309 241226 293375 241229
rect 147121 241224 277410 241226
rect -960 241090 480 241180
rect 147121 241168 147126 241224
rect 147182 241168 277410 241224
rect 147121 241166 277410 241168
rect 292806 241224 293375 241226
rect 292806 241168 293314 241224
rect 293370 241168 293375 241224
rect 292806 241166 293375 241168
rect 147121 241163 147187 241166
rect 2957 241090 3023 241093
rect -960 241088 3023 241090
rect -960 241032 2962 241088
rect 3018 241032 3023 241088
rect -960 241030 3023 241032
rect 277350 241090 277410 241166
rect 293309 241163 293375 241166
rect 301129 241090 301195 241093
rect 277350 241088 301195 241090
rect 277350 241032 301134 241088
rect 301190 241032 301195 241088
rect 277350 241030 301195 241032
rect -960 240940 480 241030
rect 2957 241027 3023 241030
rect 301129 241027 301195 241030
rect 119889 240954 119955 240957
rect 128353 240954 128419 240957
rect 119889 240952 128419 240954
rect 119889 240896 119894 240952
rect 119950 240896 128358 240952
rect 128414 240896 128419 240952
rect 119889 240894 128419 240896
rect 119889 240891 119955 240894
rect 128353 240891 128419 240894
rect 67633 240818 67699 240821
rect 121453 240818 121519 240821
rect 67633 240816 70196 240818
rect 67633 240760 67638 240816
rect 67694 240760 70196 240816
rect 67633 240758 70196 240760
rect 119876 240816 121519 240818
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 67633 240755 67699 240758
rect 121453 240755 121519 240758
rect 165521 240818 165587 240821
rect 165521 240816 200130 240818
rect 165521 240760 165526 240816
rect 165582 240760 200130 240816
rect 165521 240758 200130 240760
rect 165521 240755 165587 240758
rect 200070 240682 200130 240758
rect 298502 240756 298508 240820
rect 298572 240818 298578 240820
rect 580257 240818 580323 240821
rect 298572 240816 580323 240818
rect 298572 240760 580262 240816
rect 580318 240760 580323 240816
rect 298572 240758 580323 240760
rect 298572 240756 298578 240758
rect 580257 240755 580323 240758
rect 215293 240682 215359 240685
rect 200070 240680 215359 240682
rect 200070 240624 215298 240680
rect 215354 240624 215359 240680
rect 200070 240622 215359 240624
rect 215293 240619 215359 240622
rect 121545 240138 121611 240141
rect 119876 240136 121611 240138
rect 119876 240080 121550 240136
rect 121606 240080 121611 240136
rect 119876 240078 121611 240080
rect 121545 240075 121611 240078
rect 287697 240138 287763 240141
rect 295374 240138 295380 240140
rect 287697 240136 295380 240138
rect 287697 240080 287702 240136
rect 287758 240080 295380 240136
rect 287697 240078 295380 240080
rect 287697 240075 287763 240078
rect 295374 240076 295380 240078
rect 295444 240076 295450 240140
rect 61745 239458 61811 239461
rect 61745 239456 103530 239458
rect 61745 239400 61750 239456
rect 61806 239400 103530 239456
rect 61745 239398 103530 239400
rect 61745 239395 61811 239398
rect 103470 239322 103530 239398
rect 111149 239322 111215 239325
rect 103470 239320 111215 239322
rect 103470 239264 111154 239320
rect 111210 239264 111215 239320
rect 103470 239262 111215 239264
rect 111149 239259 111215 239262
rect 292665 239188 292731 239189
rect 292614 239124 292620 239188
rect 292684 239186 292731 239188
rect 292684 239184 292776 239186
rect 292726 239128 292776 239184
rect 292684 239126 292776 239128
rect 292684 239124 292731 239126
rect 292665 239123 292731 239124
rect 56225 238778 56291 238781
rect 74533 238778 74599 238781
rect 56225 238776 74599 238778
rect 56225 238720 56230 238776
rect 56286 238720 74538 238776
rect 74594 238720 74599 238776
rect 56225 238718 74599 238720
rect 56225 238715 56291 238718
rect 74533 238715 74599 238718
rect 109033 238778 109099 238781
rect 109953 238778 110019 238781
rect 124070 238778 124076 238780
rect 109033 238776 124076 238778
rect 109033 238720 109038 238776
rect 109094 238720 109958 238776
rect 110014 238720 124076 238776
rect 109033 238718 124076 238720
rect 109033 238715 109099 238718
rect 109953 238715 110019 238718
rect 124070 238716 124076 238718
rect 124140 238716 124146 238780
rect 167821 238778 167887 238781
rect 224033 238778 224099 238781
rect 314653 238778 314719 238781
rect 167821 238776 314719 238778
rect 167821 238720 167826 238776
rect 167882 238720 224038 238776
rect 224094 238720 314658 238776
rect 314714 238720 314719 238776
rect 167821 238718 314719 238720
rect 167821 238715 167887 238718
rect 224033 238715 224099 238718
rect 314653 238715 314719 238718
rect 57830 238580 57836 238644
rect 57900 238642 57906 238644
rect 72601 238642 72667 238645
rect 57900 238640 72667 238642
rect 57900 238584 72606 238640
rect 72662 238584 72667 238640
rect 57900 238582 72667 238584
rect 57900 238580 57906 238582
rect 72601 238579 72667 238582
rect 86125 238642 86191 238645
rect 158621 238642 158687 238645
rect 86125 238640 158687 238642
rect 86125 238584 86130 238640
rect 86186 238584 158626 238640
rect 158682 238584 158687 238640
rect 86125 238582 158687 238584
rect 86125 238579 86191 238582
rect 158621 238579 158687 238582
rect 161974 238580 161980 238644
rect 162044 238642 162050 238644
rect 582465 238642 582531 238645
rect 162044 238640 582531 238642
rect 162044 238584 582470 238640
rect 582526 238584 582531 238640
rect 162044 238582 582531 238584
rect 162044 238580 162050 238582
rect 582465 238579 582531 238582
rect 66897 238506 66963 238509
rect 117681 238506 117747 238509
rect 66897 238504 117747 238506
rect 66897 238448 66902 238504
rect 66958 238448 117686 238504
rect 117742 238448 117747 238504
rect 66897 238446 117747 238448
rect 66897 238443 66963 238446
rect 117681 238443 117747 238446
rect 158621 237418 158687 237421
rect 160737 237418 160803 237421
rect 158621 237416 160803 237418
rect 158621 237360 158626 237416
rect 158682 237360 160742 237416
rect 160798 237360 160803 237416
rect 158621 237358 160803 237360
rect 158621 237355 158687 237358
rect 160737 237355 160803 237358
rect 184197 237418 184263 237421
rect 184790 237418 184796 237420
rect 184197 237416 184796 237418
rect 184197 237360 184202 237416
rect 184258 237360 184796 237416
rect 184197 237358 184796 237360
rect 184197 237355 184263 237358
rect 184790 237356 184796 237358
rect 184860 237356 184866 237420
rect 61878 237220 61884 237284
rect 61948 237282 61954 237284
rect 163497 237282 163563 237285
rect 61948 237280 163563 237282
rect 61948 237224 163502 237280
rect 163558 237224 163563 237280
rect 61948 237222 163563 237224
rect 61948 237220 61954 237222
rect 163497 237219 163563 237222
rect 72601 237146 72667 237149
rect 120574 237146 120580 237148
rect 72601 237144 120580 237146
rect 72601 237088 72606 237144
rect 72662 237088 120580 237144
rect 72601 237086 120580 237088
rect 72601 237083 72667 237086
rect 120574 237084 120580 237086
rect 120644 237084 120650 237148
rect 114461 237010 114527 237013
rect 134374 237010 134380 237012
rect 114461 237008 134380 237010
rect 114461 236952 114466 237008
rect 114522 236952 134380 237008
rect 114461 236950 134380 236952
rect 114461 236947 114527 236950
rect 134374 236948 134380 236950
rect 134444 236948 134450 237012
rect 275277 235378 275343 235381
rect 293166 235378 293172 235380
rect 275277 235376 293172 235378
rect 275277 235320 275282 235376
rect 275338 235320 293172 235376
rect 275277 235318 293172 235320
rect 275277 235315 275343 235318
rect 293166 235316 293172 235318
rect 293236 235316 293242 235380
rect 64454 235180 64460 235244
rect 64524 235242 64530 235244
rect 314561 235242 314627 235245
rect 323025 235242 323091 235245
rect 64524 235240 323091 235242
rect 64524 235184 314566 235240
rect 314622 235184 323030 235240
rect 323086 235184 323091 235240
rect 64524 235182 323091 235184
rect 64524 235180 64530 235182
rect 314561 235179 314627 235182
rect 323025 235179 323091 235182
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 169702 231780 169708 231844
rect 169772 231842 169778 231844
rect 170765 231842 170831 231845
rect 169772 231840 170831 231842
rect 169772 231784 170770 231840
rect 170826 231784 170831 231840
rect 169772 231782 170831 231784
rect 169772 231780 169778 231782
rect 170765 231779 170831 231782
rect 179781 231844 179847 231845
rect 179781 231840 179828 231844
rect 179892 231842 179898 231844
rect 179781 231784 179786 231840
rect 179781 231780 179828 231784
rect 179892 231782 179938 231842
rect 179892 231780 179898 231782
rect 179781 231779 179847 231780
rect 122097 228986 122163 228989
rect 331254 228986 331260 228988
rect 122097 228984 331260 228986
rect 122097 228928 122102 228984
rect 122158 228928 331260 228984
rect 122097 228926 331260 228928
rect 122097 228923 122163 228926
rect 331254 228924 331260 228926
rect 331324 228924 331330 228988
rect -960 227884 480 228124
rect 328545 227762 328611 227765
rect 328678 227762 328684 227764
rect 328545 227760 328684 227762
rect 328545 227704 328550 227760
rect 328606 227704 328684 227760
rect 328545 227702 328684 227704
rect 328545 227699 328611 227702
rect 328678 227700 328684 227702
rect 328748 227700 328754 227764
rect 179086 226884 179092 226948
rect 179156 226946 179162 226948
rect 580349 226946 580415 226949
rect 179156 226944 580415 226946
rect 179156 226888 580354 226944
rect 580410 226888 580415 226944
rect 179156 226886 580415 226888
rect 179156 226884 179162 226886
rect 580349 226883 580415 226886
rect 178769 226402 178835 226405
rect 178902 226402 178908 226404
rect 178769 226400 178908 226402
rect 178769 226344 178774 226400
rect 178830 226344 178908 226400
rect 178769 226342 178908 226344
rect 178769 226339 178835 226342
rect 178902 226340 178908 226342
rect 178972 226340 178978 226404
rect 54845 225586 54911 225589
rect 256734 225586 256740 225588
rect 54845 225584 256740 225586
rect 54845 225528 54850 225584
rect 54906 225528 256740 225584
rect 54845 225526 256740 225528
rect 54845 225523 54911 225526
rect 256734 225524 256740 225526
rect 256804 225524 256810 225588
rect 161473 224226 161539 224229
rect 259494 224226 259500 224228
rect 161473 224224 259500 224226
rect 161473 224168 161478 224224
rect 161534 224168 259500 224224
rect 161473 224166 259500 224168
rect 161473 224163 161539 224166
rect 259494 224164 259500 224166
rect 259564 224164 259570 224228
rect 324313 223682 324379 223685
rect 324957 223682 325023 223685
rect 338246 223682 338252 223684
rect 324313 223680 338252 223682
rect 324313 223624 324318 223680
rect 324374 223624 324962 223680
rect 325018 223624 338252 223680
rect 324313 223622 338252 223624
rect 324313 223619 324379 223622
rect 324957 223619 325023 223622
rect 338246 223620 338252 223622
rect 338316 223620 338322 223684
rect 85481 222866 85547 222869
rect 252502 222866 252508 222868
rect 85481 222864 252508 222866
rect 85481 222808 85486 222864
rect 85542 222808 252508 222864
rect 85481 222806 252508 222808
rect 85481 222803 85547 222806
rect 252502 222804 252508 222806
rect 252572 222804 252578 222868
rect 63166 222124 63172 222188
rect 63236 222186 63242 222188
rect 262213 222186 262279 222189
rect 262857 222186 262923 222189
rect 63236 222184 262923 222186
rect 63236 222128 262218 222184
rect 262274 222128 262862 222184
rect 262918 222128 262923 222184
rect 63236 222126 262923 222128
rect 63236 222124 63242 222126
rect 262213 222123 262279 222126
rect 262857 222123 262923 222126
rect 149646 221988 149652 222052
rect 149716 222050 149722 222052
rect 336733 222050 336799 222053
rect 149716 222048 336799 222050
rect 149716 221992 336738 222048
rect 336794 221992 336799 222048
rect 149716 221990 336799 221992
rect 149716 221988 149722 221990
rect 336733 221987 336799 221990
rect 329833 220828 329899 220829
rect 166390 220764 166396 220828
rect 166460 220826 166466 220828
rect 329782 220826 329788 220828
rect 166460 220766 329788 220826
rect 329852 220824 329899 220828
rect 329894 220768 329899 220824
rect 166460 220764 166466 220766
rect 329782 220764 329788 220766
rect 329852 220764 329899 220768
rect 329833 220763 329899 220764
rect 327073 219332 327139 219333
rect 327022 219268 327028 219332
rect 327092 219330 327139 219332
rect 327092 219328 327184 219330
rect 327134 219272 327184 219328
rect 327092 219270 327184 219272
rect 327092 219268 327139 219270
rect 327073 219267 327139 219268
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 130326 213148 130332 213212
rect 130396 213210 130402 213212
rect 336774 213210 336780 213212
rect 130396 213150 336780 213210
rect 130396 213148 130402 213150
rect 336774 213148 336780 213150
rect 336844 213148 336850 213212
rect 119838 210292 119844 210356
rect 119908 210354 119914 210356
rect 325693 210354 325759 210357
rect 119908 210352 325759 210354
rect 119908 210296 325698 210352
rect 325754 210296 325759 210352
rect 119908 210294 325759 210296
rect 119908 210292 119914 210294
rect 325693 210291 325759 210294
rect 579889 205730 579955 205733
rect 583520 205730 584960 205820
rect 579889 205728 584960 205730
rect 579889 205672 579894 205728
rect 579950 205672 584960 205728
rect 579889 205670 584960 205672
rect 579889 205667 579955 205670
rect 583520 205580 584960 205670
rect 129181 204914 129247 204917
rect 265014 204914 265020 204916
rect 129181 204912 265020 204914
rect 129181 204856 129186 204912
rect 129242 204856 265020 204912
rect 129181 204854 265020 204856
rect 129181 204851 129247 204854
rect 265014 204852 265020 204854
rect 265084 204852 265090 204916
rect 57697 202330 57763 202333
rect 260966 202330 260972 202332
rect 57697 202328 260972 202330
rect 57697 202272 57702 202328
rect 57758 202272 260972 202328
rect 57697 202270 260972 202272
rect 57697 202267 57763 202270
rect 260966 202268 260972 202270
rect 261036 202268 261042 202332
rect 128854 202132 128860 202196
rect 128924 202194 128930 202196
rect 339493 202194 339559 202197
rect 128924 202192 339559 202194
rect 128924 202136 339498 202192
rect 339554 202136 339559 202192
rect 128924 202134 339559 202136
rect 128924 202132 128930 202134
rect 339493 202131 339559 202134
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 52177 200834 52243 200837
rect 266302 200834 266308 200836
rect 52177 200832 266308 200834
rect 52177 200776 52182 200832
rect 52238 200776 266308 200832
rect 52177 200774 266308 200776
rect 52177 200771 52243 200774
rect 266302 200772 266308 200774
rect 266372 200772 266378 200836
rect 64638 200636 64644 200700
rect 64708 200698 64714 200700
rect 342437 200698 342503 200701
rect 64708 200696 342503 200698
rect 64708 200640 342442 200696
rect 342498 200640 342503 200696
rect 64708 200638 342503 200640
rect 64708 200636 64714 200638
rect 342437 200635 342503 200638
rect 327574 196692 327580 196756
rect 327644 196754 327650 196756
rect 336733 196754 336799 196757
rect 327644 196752 336799 196754
rect 327644 196696 336738 196752
rect 336794 196696 336799 196752
rect 327644 196694 336799 196696
rect 327644 196692 327650 196694
rect 336733 196691 336799 196694
rect 138606 196556 138612 196620
rect 138676 196618 138682 196620
rect 345054 196618 345060 196620
rect 138676 196558 345060 196618
rect 138676 196556 138682 196558
rect 345054 196556 345060 196558
rect 345124 196556 345130 196620
rect 117957 195258 118023 195261
rect 335670 195258 335676 195260
rect 117957 195256 335676 195258
rect 117957 195200 117962 195256
rect 118018 195200 335676 195256
rect 117957 195198 335676 195200
rect 117957 195195 118023 195198
rect 335670 195196 335676 195198
rect 335740 195196 335746 195260
rect 149881 194034 149947 194037
rect 257838 194034 257844 194036
rect 149881 194032 257844 194034
rect 149881 193976 149886 194032
rect 149942 193976 257844 194032
rect 149881 193974 257844 193976
rect 149881 193971 149947 193974
rect 257838 193972 257844 193974
rect 257908 193972 257914 194036
rect 67398 193836 67404 193900
rect 67468 193898 67474 193900
rect 324405 193898 324471 193901
rect 67468 193896 324471 193898
rect 67468 193840 324410 193896
rect 324466 193840 324471 193896
rect 67468 193838 324471 193840
rect 67468 193836 67474 193838
rect 324405 193835 324471 193838
rect 162301 192538 162367 192541
rect 263726 192538 263732 192540
rect 162301 192536 263732 192538
rect 162301 192480 162306 192536
rect 162362 192480 263732 192536
rect 162301 192478 263732 192480
rect 162301 192475 162367 192478
rect 263726 192476 263732 192478
rect 263796 192476 263802 192540
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect 224953 191178 225019 191181
rect 269614 191178 269620 191180
rect 224953 191176 269620 191178
rect 224953 191120 224958 191176
rect 225014 191120 269620 191176
rect 224953 191118 269620 191120
rect 224953 191115 225019 191118
rect 269614 191116 269620 191118
rect 269684 191116 269690 191180
rect 152641 191042 152707 191045
rect 260782 191042 260788 191044
rect 152641 191040 260788 191042
rect 152641 190984 152646 191040
rect 152702 190984 260788 191040
rect 152641 190982 260788 190984
rect 152641 190979 152707 190982
rect 260782 190980 260788 190982
rect 260852 190980 260858 191044
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 229093 188594 229159 188597
rect 271086 188594 271092 188596
rect 229093 188592 271092 188594
rect 229093 188536 229098 188592
rect 229154 188536 271092 188592
rect 229093 188534 271092 188536
rect 229093 188531 229159 188534
rect 271086 188532 271092 188534
rect 271156 188532 271162 188596
rect 142797 188458 142863 188461
rect 263542 188458 263548 188460
rect 142797 188456 263548 188458
rect 142797 188400 142802 188456
rect 142858 188400 263548 188456
rect 142797 188398 263548 188400
rect 142797 188395 142863 188398
rect 263542 188396 263548 188398
rect 263612 188396 263618 188460
rect 148174 188260 148180 188324
rect 148244 188322 148250 188324
rect 339677 188322 339743 188325
rect 148244 188320 339743 188322
rect 148244 188264 339682 188320
rect 339738 188264 339743 188320
rect 148244 188262 339743 188264
rect 148244 188260 148250 188262
rect 339677 188259 339743 188262
rect 151077 186962 151143 186965
rect 318006 186962 318012 186964
rect 151077 186960 318012 186962
rect 151077 186904 151082 186960
rect 151138 186904 318012 186960
rect 151077 186902 318012 186904
rect 151077 186899 151143 186902
rect 318006 186900 318012 186902
rect 318076 186900 318082 186964
rect 250437 186418 250503 186421
rect 255446 186418 255452 186420
rect 250437 186416 255452 186418
rect 250437 186360 250442 186416
rect 250498 186360 255452 186416
rect 250437 186358 255452 186360
rect 250437 186355 250503 186358
rect 255446 186356 255452 186358
rect 255516 186356 255522 186420
rect 80697 185602 80763 185605
rect 320214 185602 320220 185604
rect 80697 185600 320220 185602
rect 80697 185544 80702 185600
rect 80758 185544 320220 185600
rect 80697 185542 320220 185544
rect 80697 185539 80763 185542
rect 320214 185540 320220 185542
rect 320284 185540 320290 185604
rect 153694 184180 153700 184244
rect 153764 184242 153770 184244
rect 336917 184242 336983 184245
rect 153764 184240 336983 184242
rect 153764 184184 336922 184240
rect 336978 184184 336983 184240
rect 153764 184182 336983 184184
rect 153764 184180 153770 184182
rect 336917 184179 336983 184182
rect 151169 182882 151235 182885
rect 265198 182882 265204 182884
rect 151169 182880 265204 182882
rect 151169 182824 151174 182880
rect 151230 182824 265204 182880
rect 151169 182822 265204 182824
rect 151169 182819 151235 182822
rect 265198 182820 265204 182822
rect 265268 182820 265274 182884
rect 114001 182202 114067 182205
rect 166390 182202 166396 182204
rect 114001 182200 166396 182202
rect 114001 182144 114006 182200
rect 114062 182144 166396 182200
rect 114001 182142 166396 182144
rect 114001 182139 114067 182142
rect 166390 182140 166396 182142
rect 166460 182140 166466 182204
rect 130377 181658 130443 181661
rect 169702 181658 169708 181660
rect 130377 181656 169708 181658
rect 130377 181600 130382 181656
rect 130438 181600 169708 181656
rect 130377 181598 169708 181600
rect 130377 181595 130443 181598
rect 169702 181596 169708 181598
rect 169772 181596 169778 181660
rect 164877 181522 164943 181525
rect 255262 181522 255268 181524
rect 164877 181520 255268 181522
rect 164877 181464 164882 181520
rect 164938 181464 255268 181520
rect 164877 181462 255268 181464
rect 164877 181459 164943 181462
rect 255262 181460 255268 181462
rect 255332 181460 255338 181524
rect 68921 181386 68987 181389
rect 322054 181386 322060 181388
rect 68921 181384 322060 181386
rect 68921 181328 68926 181384
rect 68982 181328 322060 181384
rect 68921 181326 322060 181328
rect 68921 181323 68987 181326
rect 322054 181324 322060 181326
rect 322124 181324 322130 181388
rect 166206 180100 166212 180164
rect 166276 180162 166282 180164
rect 335670 180162 335676 180164
rect 166276 180102 335676 180162
rect 166276 180100 166282 180102
rect 335670 180100 335676 180102
rect 335740 180100 335746 180164
rect 160686 179964 160692 180028
rect 160756 180026 160762 180028
rect 343909 180026 343975 180029
rect 160756 180024 343975 180026
rect 160756 179968 343914 180024
rect 343970 179968 343975 180024
rect 160756 179966 343975 179968
rect 160756 179964 160762 179966
rect 343909 179963 343975 179966
rect 346301 179348 346367 179349
rect 346301 179346 346348 179348
rect 346256 179344 346348 179346
rect 346256 179288 346306 179344
rect 346256 179286 346348 179288
rect 346301 179284 346348 179286
rect 346412 179284 346418 179348
rect 346301 179283 346367 179284
rect 342294 179148 342300 179212
rect 342364 179210 342370 179212
rect 342621 179210 342687 179213
rect 342364 179208 342687 179210
rect 342364 179152 342626 179208
rect 342682 179152 342687 179208
rect 342364 179150 342687 179152
rect 342364 179148 342370 179150
rect 342621 179147 342687 179150
rect 580257 179210 580323 179213
rect 583520 179210 584960 179300
rect 580257 179208 584960 179210
rect 580257 179152 580262 179208
rect 580318 179152 584960 179208
rect 580257 179150 584960 179152
rect 580257 179147 580323 179150
rect 583520 179060 584960 179150
rect 231117 178938 231183 178941
rect 249006 178938 249012 178940
rect 231117 178936 249012 178938
rect 231117 178880 231122 178936
rect 231178 178880 249012 178936
rect 231117 178878 249012 178880
rect 231117 178875 231183 178878
rect 249006 178876 249012 178878
rect 249076 178876 249082 178940
rect 239397 178802 239463 178805
rect 259678 178802 259684 178804
rect 239397 178800 259684 178802
rect 239397 178744 239402 178800
rect 239458 178744 259684 178800
rect 239397 178742 259684 178744
rect 239397 178739 239463 178742
rect 259678 178740 259684 178742
rect 259748 178740 259754 178804
rect 162117 178666 162183 178669
rect 256918 178666 256924 178668
rect 162117 178664 256924 178666
rect 162117 178608 162122 178664
rect 162178 178608 256924 178664
rect 162117 178606 256924 178608
rect 162117 178603 162183 178606
rect 256918 178604 256924 178606
rect 256988 178604 256994 178668
rect 283649 178666 283715 178669
rect 332726 178666 332732 178668
rect 283649 178664 332732 178666
rect 283649 178608 283654 178664
rect 283710 178608 332732 178664
rect 283649 178606 332732 178608
rect 283649 178603 283715 178606
rect 332726 178604 332732 178606
rect 332796 178604 332802 178668
rect 110638 178196 110644 178260
rect 110708 178258 110714 178260
rect 167678 178258 167684 178260
rect 110708 178198 167684 178258
rect 110708 178196 110714 178198
rect 167678 178196 167684 178198
rect 167748 178196 167754 178260
rect 166206 178122 166212 178124
rect 97030 178062 166212 178122
rect 97030 177988 97090 178062
rect 166206 178060 166212 178062
rect 166276 178060 166282 178124
rect 97022 177924 97028 177988
rect 97092 177924 97098 177988
rect 99414 177516 99420 177580
rect 99484 177578 99490 177580
rect 100661 177578 100727 177581
rect 102041 177580 102107 177581
rect 101990 177578 101996 177580
rect 99484 177576 100727 177578
rect 99484 177520 100666 177576
rect 100722 177520 100727 177576
rect 99484 177518 100727 177520
rect 101950 177518 101996 177578
rect 102060 177576 102107 177580
rect 102102 177520 102107 177576
rect 99484 177516 99490 177518
rect 100661 177515 100727 177518
rect 101990 177516 101996 177518
rect 102060 177516 102107 177520
rect 104566 177516 104572 177580
rect 104636 177578 104642 177580
rect 104801 177578 104867 177581
rect 104636 177576 104867 177578
rect 104636 177520 104806 177576
rect 104862 177520 104867 177576
rect 104636 177518 104867 177520
rect 104636 177516 104642 177518
rect 102041 177515 102107 177516
rect 104801 177515 104867 177518
rect 106038 177516 106044 177580
rect 106108 177578 106114 177580
rect 106181 177578 106247 177581
rect 106108 177576 106247 177578
rect 106108 177520 106186 177576
rect 106242 177520 106247 177576
rect 106108 177518 106247 177520
rect 106108 177516 106114 177518
rect 106181 177515 106247 177518
rect 113214 177516 113220 177580
rect 113284 177578 113290 177580
rect 114001 177578 114067 177581
rect 118417 177580 118483 177581
rect 118366 177578 118372 177580
rect 113284 177576 114067 177578
rect 113284 177520 114006 177576
rect 114062 177520 114067 177576
rect 113284 177518 114067 177520
rect 118326 177518 118372 177578
rect 118436 177576 118483 177580
rect 118478 177520 118483 177576
rect 113284 177516 113290 177518
rect 114001 177515 114067 177518
rect 118366 177516 118372 177518
rect 118436 177516 118483 177520
rect 121862 177516 121868 177580
rect 121932 177578 121938 177580
rect 122005 177578 122071 177581
rect 121932 177576 122071 177578
rect 121932 177520 122010 177576
rect 122066 177520 122071 177576
rect 121932 177518 122071 177520
rect 121932 177516 121938 177518
rect 118417 177515 118483 177516
rect 122005 177515 122071 177518
rect 124438 177516 124444 177580
rect 124508 177578 124514 177580
rect 125501 177578 125567 177581
rect 124508 177576 125567 177578
rect 124508 177520 125506 177576
rect 125562 177520 125567 177576
rect 124508 177518 125567 177520
rect 124508 177516 124514 177518
rect 125501 177515 125567 177518
rect 131982 177516 131988 177580
rect 132052 177578 132058 177580
rect 132401 177578 132467 177581
rect 132052 177576 132467 177578
rect 132052 177520 132406 177576
rect 132462 177520 132467 177576
rect 132052 177518 132467 177520
rect 132052 177516 132058 177518
rect 132401 177515 132467 177518
rect 133086 177516 133092 177580
rect 133156 177578 133162 177580
rect 133597 177578 133663 177581
rect 133156 177576 133663 177578
rect 133156 177520 133602 177576
rect 133658 177520 133663 177576
rect 133156 177518 133663 177520
rect 133156 177516 133162 177518
rect 133597 177515 133663 177518
rect 248505 177578 248571 177581
rect 249190 177578 249196 177580
rect 248505 177576 249196 177578
rect 248505 177520 248510 177576
rect 248566 177520 249196 177576
rect 248505 177518 249196 177520
rect 248505 177515 248571 177518
rect 249190 177516 249196 177518
rect 249260 177516 249266 177580
rect 318006 177516 318012 177580
rect 318076 177578 318082 177580
rect 325969 177578 326035 177581
rect 318076 177576 326035 177578
rect 318076 177520 325974 177576
rect 326030 177520 326035 177576
rect 318076 177518 326035 177520
rect 318076 177516 318082 177518
rect 325969 177515 326035 177518
rect 318149 177442 318215 177445
rect 334014 177442 334020 177444
rect 318149 177440 334020 177442
rect 318149 177384 318154 177440
rect 318210 177384 334020 177440
rect 318149 177382 334020 177384
rect 318149 177379 318215 177382
rect 334014 177380 334020 177382
rect 334084 177380 334090 177444
rect 1301 177306 1367 177309
rect 52545 177308 52611 177309
rect 52494 177306 52500 177308
rect 1301 177304 52500 177306
rect 52564 177306 52611 177308
rect 166901 177306 166967 177309
rect 206277 177306 206343 177309
rect 52564 177304 52692 177306
rect 1301 177248 1306 177304
rect 1362 177248 52500 177304
rect 52606 177248 52692 177304
rect 1301 177246 52500 177248
rect 1301 177243 1367 177246
rect 52494 177244 52500 177246
rect 52564 177246 52692 177248
rect 166901 177304 206343 177306
rect 166901 177248 166906 177304
rect 166962 177248 206282 177304
rect 206338 177248 206343 177304
rect 166901 177246 206343 177248
rect 52564 177244 52611 177246
rect 52545 177243 52611 177244
rect 166901 177243 166967 177246
rect 206277 177243 206343 177246
rect 246389 177306 246455 177309
rect 254117 177306 254183 177309
rect 246389 177304 254183 177306
rect 246389 177248 246394 177304
rect 246450 177248 254122 177304
rect 254178 177248 254183 177304
rect 246389 177246 254183 177248
rect 246389 177243 246455 177246
rect 254117 177243 254183 177246
rect 307109 177306 307175 177309
rect 336958 177306 336964 177308
rect 307109 177304 336964 177306
rect 307109 177248 307114 177304
rect 307170 177248 336964 177304
rect 307109 177246 336964 177248
rect 307109 177243 307175 177246
rect 336958 177244 336964 177246
rect 337028 177244 337034 177308
rect 114134 176972 114140 177036
rect 114204 177034 114210 177036
rect 114277 177034 114343 177037
rect 114204 177032 114343 177034
rect 114204 176976 114282 177032
rect 114338 176976 114343 177032
rect 114204 176974 114343 176976
rect 114204 176972 114210 176974
rect 114277 176971 114343 176974
rect 120758 176972 120764 177036
rect 120828 177034 120834 177036
rect 120993 177034 121059 177037
rect 123017 177036 123083 177037
rect 122966 177034 122972 177036
rect 120828 177032 121059 177034
rect 120828 176976 120998 177032
rect 121054 176976 121059 177032
rect 120828 176974 121059 176976
rect 122926 176974 122972 177034
rect 123036 177032 123083 177036
rect 123078 176976 123083 177032
rect 120828 176972 120834 176974
rect 120993 176971 121059 176974
rect 122966 176972 122972 176974
rect 123036 176972 123083 176976
rect 123017 176971 123083 176972
rect 103278 176836 103284 176900
rect 103348 176898 103354 176900
rect 167494 176898 167500 176900
rect 103348 176838 167500 176898
rect 103348 176836 103354 176838
rect 167494 176836 167500 176838
rect 167564 176836 167570 176900
rect 107009 176764 107075 176765
rect 108113 176764 108179 176765
rect 106958 176762 106964 176764
rect 106918 176702 106964 176762
rect 107028 176760 107075 176764
rect 108062 176762 108068 176764
rect 107070 176704 107075 176760
rect 106958 176700 106964 176702
rect 107028 176700 107075 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 109953 176762 110019 176765
rect 109604 176760 110019 176762
rect 109604 176704 109958 176760
rect 110014 176704 110019 176760
rect 109604 176702 110019 176704
rect 109604 176700 109610 176702
rect 107009 176699 107075 176700
rect 108113 176699 108179 176700
rect 109953 176699 110019 176702
rect 112110 176700 112116 176764
rect 112180 176762 112186 176764
rect 112437 176762 112503 176765
rect 125777 176764 125843 176765
rect 127065 176764 127131 176765
rect 125726 176762 125732 176764
rect 112180 176760 112503 176762
rect 112180 176704 112442 176760
rect 112498 176704 112503 176760
rect 112180 176702 112503 176704
rect 125686 176702 125732 176762
rect 125796 176760 125843 176764
rect 127014 176762 127020 176764
rect 125838 176704 125843 176760
rect 112180 176700 112186 176702
rect 112437 176699 112503 176702
rect 125726 176700 125732 176702
rect 125796 176700 125843 176704
rect 126974 176702 127020 176762
rect 127084 176760 127131 176764
rect 128169 176762 128235 176765
rect 130745 176764 130811 176765
rect 134425 176764 134491 176765
rect 135713 176764 135779 176765
rect 148225 176764 148291 176765
rect 130694 176762 130700 176764
rect 127126 176704 127131 176760
rect 127014 176700 127020 176702
rect 127084 176700 127131 176704
rect 125777 176699 125843 176700
rect 127065 176699 127131 176700
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 130654 176702 130700 176762
rect 130764 176760 130811 176764
rect 134374 176762 134380 176764
rect 130806 176704 130811 176760
rect 130694 176700 130700 176702
rect 130764 176700 130811 176704
rect 134334 176702 134380 176762
rect 134444 176760 134491 176764
rect 135662 176762 135668 176764
rect 134486 176704 134491 176760
rect 134374 176700 134380 176702
rect 134444 176700 134491 176704
rect 135622 176702 135668 176762
rect 135732 176760 135779 176764
rect 148174 176762 148180 176764
rect 135774 176704 135779 176760
rect 135662 176700 135668 176702
rect 135732 176700 135779 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 159909 176762 159975 176765
rect 158916 176760 159975 176762
rect 158916 176704 159914 176760
rect 159970 176704 159975 176760
rect 158916 176702 159975 176704
rect 158916 176700 158922 176702
rect 130745 176699 130811 176700
rect 134425 176699 134491 176700
rect 135713 176699 135779 176700
rect 148225 176699 148291 176700
rect 159909 176699 159975 176702
rect 128126 176492 128186 176699
rect 162393 176626 162459 176629
rect 166533 176626 166599 176629
rect 162393 176624 166599 176626
rect 162393 176568 162398 176624
rect 162454 176568 166538 176624
rect 166594 176568 166599 176624
rect 162393 176566 166599 176568
rect 162393 176563 162459 176566
rect 166533 176563 166599 176566
rect 318425 176626 318491 176629
rect 323025 176626 323091 176629
rect 318425 176624 323091 176626
rect 318425 176568 318430 176624
rect 318486 176568 323030 176624
rect 323086 176568 323091 176624
rect 318425 176566 323091 176568
rect 318425 176563 318491 176566
rect 323025 176563 323091 176566
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 318241 176218 318307 176221
rect 321502 176218 321508 176220
rect 318241 176216 321508 176218
rect 318241 176160 318246 176216
rect 318302 176160 321508 176216
rect 318241 176158 321508 176160
rect 318241 176155 318307 176158
rect 321502 176156 321508 176158
rect 321572 176156 321578 176220
rect 247677 176082 247743 176085
rect 262254 176082 262260 176084
rect 247677 176080 262260 176082
rect -960 175796 480 176036
rect 247677 176024 247682 176080
rect 247738 176024 262260 176080
rect 247677 176022 262260 176024
rect 247677 176019 247743 176022
rect 262254 176020 262260 176022
rect 262324 176020 262330 176084
rect 321461 176082 321527 176085
rect 321461 176080 321570 176082
rect 321461 176024 321466 176080
rect 321522 176024 321570 176080
rect 321461 176019 321570 176024
rect 152549 175946 152615 175949
rect 249149 175946 249215 175949
rect 152549 175944 249215 175946
rect 152549 175888 152554 175944
rect 152610 175888 249154 175944
rect 249210 175888 249215 175944
rect 152549 175886 249215 175888
rect 152549 175883 152615 175886
rect 249149 175883 249215 175886
rect 248045 175810 248111 175813
rect 248045 175808 248338 175810
rect 248045 175752 248050 175808
rect 248106 175752 248338 175808
rect 248045 175750 248338 175752
rect 248045 175747 248111 175750
rect 213913 175674 213979 175677
rect 213913 175672 217212 175674
rect 213913 175616 213918 175672
rect 213974 175616 217212 175672
rect 248278 175644 248338 175750
rect 307017 175676 307083 175677
rect 306966 175674 306972 175676
rect 213913 175614 217212 175616
rect 306890 175614 306972 175674
rect 307036 175674 307083 175676
rect 307036 175672 310132 175674
rect 307078 175616 310132 175672
rect 213913 175611 213979 175614
rect 306966 175612 306972 175614
rect 307036 175614 310132 175616
rect 307036 175612 307083 175614
rect 307017 175611 307083 175612
rect 321510 175508 321570 176019
rect 98361 175404 98427 175405
rect 100753 175404 100819 175405
rect 116945 175404 117011 175405
rect 129457 175404 129523 175405
rect 98310 175402 98316 175404
rect 98270 175342 98316 175402
rect 98380 175400 98427 175404
rect 100702 175402 100708 175404
rect 98422 175344 98427 175400
rect 98310 175340 98316 175342
rect 98380 175340 98427 175344
rect 100662 175342 100708 175402
rect 100772 175400 100819 175404
rect 116894 175402 116900 175404
rect 100814 175344 100819 175400
rect 100702 175340 100708 175342
rect 100772 175340 100819 175344
rect 116854 175342 116900 175402
rect 116964 175400 117011 175404
rect 129406 175402 129412 175404
rect 117006 175344 117011 175400
rect 116894 175340 116900 175342
rect 116964 175340 117011 175344
rect 129366 175342 129412 175402
rect 129476 175400 129523 175404
rect 129518 175344 129523 175400
rect 129406 175340 129412 175342
rect 129476 175340 129523 175344
rect 98361 175339 98427 175340
rect 100753 175339 100819 175340
rect 116945 175339 117011 175340
rect 129457 175339 129523 175340
rect 249333 175266 249399 175269
rect 248860 175264 249399 175266
rect 248860 175208 249338 175264
rect 249394 175208 249399 175264
rect 248860 175206 249399 175208
rect 249333 175203 249399 175206
rect 307569 175266 307635 175269
rect 307569 175264 310132 175266
rect 307569 175208 307574 175264
rect 307630 175208 310132 175264
rect 307569 175206 310132 175208
rect 307569 175203 307635 175206
rect 115749 174996 115815 174997
rect 119429 174996 119495 174997
rect 115720 174994 115726 174996
rect 115658 174934 115726 174994
rect 115790 174992 115815 174996
rect 119392 174994 119398 174996
rect 115810 174936 115815 174992
rect 115720 174932 115726 174934
rect 115790 174932 115815 174936
rect 119338 174934 119398 174994
rect 119462 174992 119495 174996
rect 119490 174936 119495 174992
rect 119392 174932 119398 174934
rect 119462 174932 119495 174936
rect 115749 174931 115815 174932
rect 119429 174931 119495 174932
rect 213913 174994 213979 174997
rect 213913 174992 217212 174994
rect 213913 174936 213918 174992
rect 213974 174936 217212 174992
rect 213913 174934 217212 174936
rect 213913 174931 213979 174934
rect 307017 174858 307083 174861
rect 307017 174856 310132 174858
rect 307017 174800 307022 174856
rect 307078 174800 310132 174856
rect 307017 174798 310132 174800
rect 307017 174795 307083 174798
rect 249149 174722 249215 174725
rect 324497 174722 324563 174725
rect 248860 174720 249215 174722
rect 248860 174664 249154 174720
rect 249210 174664 249215 174720
rect 248860 174662 249215 174664
rect 321908 174720 324563 174722
rect 321908 174664 324502 174720
rect 324558 174664 324563 174720
rect 321908 174662 324563 174664
rect 249149 174659 249215 174662
rect 324497 174659 324563 174662
rect 307293 174450 307359 174453
rect 321737 174450 321803 174453
rect 307293 174448 310132 174450
rect 307293 174392 307298 174448
rect 307354 174392 310132 174448
rect 307293 174390 310132 174392
rect 321694 174448 321803 174450
rect 321694 174392 321742 174448
rect 321798 174392 321803 174448
rect 307293 174387 307359 174390
rect 321694 174387 321803 174392
rect 214005 174314 214071 174317
rect 249190 174314 249196 174316
rect 214005 174312 217212 174314
rect 214005 174256 214010 174312
rect 214066 174256 217212 174312
rect 214005 174254 217212 174256
rect 248860 174254 249196 174314
rect 214005 174251 214071 174254
rect 249190 174252 249196 174254
rect 249260 174252 249266 174316
rect 307661 174042 307727 174045
rect 307661 174040 310132 174042
rect 307661 173984 307666 174040
rect 307722 173984 310132 174040
rect 321694 174012 321754 174387
rect 307661 173982 310132 173984
rect 307661 173979 307727 173982
rect 261017 173908 261083 173909
rect 260966 173906 260972 173908
rect 260926 173846 260972 173906
rect 261036 173904 261083 173908
rect 261078 173848 261083 173904
rect 260966 173844 260972 173846
rect 261036 173844 261083 173848
rect 261017 173843 261083 173844
rect 252461 173770 252527 173773
rect 248860 173768 252527 173770
rect 248860 173712 252466 173768
rect 252522 173712 252527 173768
rect 248860 173710 252527 173712
rect 252461 173707 252527 173710
rect 213913 173634 213979 173637
rect 307569 173634 307635 173637
rect 213913 173632 217212 173634
rect 213913 173576 213918 173632
rect 213974 173576 217212 173632
rect 213913 173574 217212 173576
rect 307569 173632 310132 173634
rect 307569 173576 307574 173632
rect 307630 173576 310132 173632
rect 307569 173574 310132 173576
rect 213913 173571 213979 173574
rect 307569 173571 307635 173574
rect 249374 173362 249380 173364
rect 248860 173302 249380 173362
rect 249374 173300 249380 173302
rect 249444 173300 249450 173364
rect 307293 173226 307359 173229
rect 323025 173226 323091 173229
rect 307293 173224 310132 173226
rect 307293 173168 307298 173224
rect 307354 173168 310132 173224
rect 307293 173166 310132 173168
rect 321908 173224 323091 173226
rect 321908 173168 323030 173224
rect 323086 173168 323091 173224
rect 321908 173166 323091 173168
rect 307293 173163 307359 173166
rect 323025 173163 323091 173166
rect 214005 172954 214071 172957
rect 214005 172952 217212 172954
rect 214005 172896 214010 172952
rect 214066 172896 217212 172952
rect 214005 172894 217212 172896
rect 214005 172891 214071 172894
rect 251725 172818 251791 172821
rect 248860 172816 251791 172818
rect 248860 172760 251730 172816
rect 251786 172760 251791 172816
rect 248860 172758 251791 172760
rect 251725 172755 251791 172758
rect 307661 172682 307727 172685
rect 321829 172682 321895 172685
rect 307661 172680 310132 172682
rect 307661 172624 307666 172680
rect 307722 172624 310132 172680
rect 307661 172622 310132 172624
rect 321829 172680 321938 172682
rect 321829 172624 321834 172680
rect 321890 172624 321938 172680
rect 307661 172619 307727 172622
rect 321829 172619 321938 172624
rect 252461 172410 252527 172413
rect 248860 172408 252527 172410
rect 248860 172352 252466 172408
rect 252522 172352 252527 172408
rect 321878 172380 321938 172619
rect 248860 172350 252527 172352
rect 252461 172347 252527 172350
rect 213913 172274 213979 172277
rect 306925 172274 306991 172277
rect 213913 172272 217212 172274
rect 213913 172216 213918 172272
rect 213974 172216 217212 172272
rect 213913 172214 217212 172216
rect 306925 172272 310132 172274
rect 306925 172216 306930 172272
rect 306986 172216 310132 172272
rect 306925 172214 310132 172216
rect 213913 172211 213979 172214
rect 306925 172211 306991 172214
rect 321502 172076 321508 172140
rect 321572 172076 321578 172140
rect 252553 171866 252619 171869
rect 248860 171864 252619 171866
rect 248860 171808 252558 171864
rect 252614 171808 252619 171864
rect 248860 171806 252619 171808
rect 252553 171803 252619 171806
rect 307477 171866 307543 171869
rect 307477 171864 310132 171866
rect 307477 171808 307482 171864
rect 307538 171808 310132 171864
rect 307477 171806 310132 171808
rect 307477 171803 307543 171806
rect 321510 171700 321570 172076
rect 167913 171594 167979 171597
rect 164694 171592 167979 171594
rect 164694 171536 167918 171592
rect 167974 171536 167979 171592
rect 164694 171534 167979 171536
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 167913 171531 167979 171534
rect 214097 171594 214163 171597
rect 214097 171592 217212 171594
rect 214097 171536 214102 171592
rect 214158 171536 217212 171592
rect 214097 171534 217212 171536
rect 214097 171531 214163 171534
rect 252369 171458 252435 171461
rect 248860 171456 252435 171458
rect 248860 171400 252374 171456
rect 252430 171400 252435 171456
rect 248860 171398 252435 171400
rect 252369 171395 252435 171398
rect 261334 171396 261340 171460
rect 261404 171458 261410 171460
rect 261404 171398 310132 171458
rect 261404 171396 261410 171398
rect 213913 171050 213979 171053
rect 307385 171050 307451 171053
rect 213913 171048 217212 171050
rect 213913 170992 213918 171048
rect 213974 170992 217212 171048
rect 213913 170990 217212 170992
rect 307385 171048 310132 171050
rect 307385 170992 307390 171048
rect 307446 170992 310132 171048
rect 307385 170990 310132 170992
rect 213913 170987 213979 170990
rect 307385 170987 307451 170990
rect 265198 170914 265204 170916
rect 248860 170854 265204 170914
rect 265198 170852 265204 170854
rect 265268 170852 265274 170916
rect 324313 170914 324379 170917
rect 321908 170912 324379 170914
rect 321908 170856 324318 170912
rect 324374 170856 324379 170912
rect 321908 170854 324379 170856
rect 324313 170851 324379 170854
rect 307477 170642 307543 170645
rect 307477 170640 310132 170642
rect 307477 170584 307482 170640
rect 307538 170584 310132 170640
rect 307477 170582 310132 170584
rect 307477 170579 307543 170582
rect 251541 170506 251607 170509
rect 248860 170504 251607 170506
rect 248860 170448 251546 170504
rect 251602 170448 251607 170504
rect 248860 170446 251607 170448
rect 251541 170443 251607 170446
rect 214005 170370 214071 170373
rect 321277 170370 321343 170373
rect 214005 170368 217212 170370
rect 214005 170312 214010 170368
rect 214066 170312 217212 170368
rect 214005 170310 217212 170312
rect 321277 170368 321386 170370
rect 321277 170312 321282 170368
rect 321338 170312 321386 170368
rect 214005 170307 214071 170310
rect 321277 170307 321386 170312
rect 307661 170234 307727 170237
rect 307661 170232 310132 170234
rect 307661 170176 307666 170232
rect 307722 170176 310132 170232
rect 307661 170174 310132 170176
rect 307661 170171 307727 170174
rect 252277 170098 252343 170101
rect 248860 170096 252343 170098
rect 248860 170040 252282 170096
rect 252338 170040 252343 170096
rect 321326 170068 321386 170307
rect 248860 170038 252343 170040
rect 252277 170035 252343 170038
rect 256785 169828 256851 169829
rect 256734 169826 256740 169828
rect 256694 169766 256740 169826
rect 256804 169824 256851 169828
rect 256846 169768 256851 169824
rect 256734 169764 256740 169766
rect 256804 169764 256851 169768
rect 256785 169763 256851 169764
rect 307293 169826 307359 169829
rect 307293 169824 310132 169826
rect 307293 169768 307298 169824
rect 307354 169768 310132 169824
rect 307293 169766 310132 169768
rect 307293 169763 307359 169766
rect 321318 169764 321324 169828
rect 321388 169826 321394 169828
rect 321388 169766 321570 169826
rect 321388 169764 321394 169766
rect 214925 169690 214991 169693
rect 214925 169688 217212 169690
rect 214925 169632 214930 169688
rect 214986 169632 217212 169688
rect 214925 169630 217212 169632
rect 214925 169627 214991 169630
rect 249977 169554 250043 169557
rect 248860 169552 250043 169554
rect 248860 169496 249982 169552
rect 250038 169496 250043 169552
rect 248860 169494 250043 169496
rect 249977 169491 250043 169494
rect 321510 169388 321570 169766
rect 307569 169282 307635 169285
rect 307569 169280 310132 169282
rect 307569 169224 307574 169280
rect 307630 169224 310132 169280
rect 307569 169222 310132 169224
rect 307569 169219 307635 169222
rect 249149 169146 249215 169149
rect 248860 169144 249215 169146
rect 248860 169088 249154 169144
rect 249210 169088 249215 169144
rect 248860 169086 249215 169088
rect 249149 169083 249215 169086
rect 213913 169010 213979 169013
rect 213913 169008 217212 169010
rect 213913 168952 213918 169008
rect 213974 168952 217212 169008
rect 213913 168950 217212 168952
rect 213913 168947 213979 168950
rect 307661 168874 307727 168877
rect 307661 168872 310132 168874
rect 307661 168816 307666 168872
rect 307722 168816 310132 168872
rect 307661 168814 310132 168816
rect 307661 168811 307727 168814
rect 252185 168602 252251 168605
rect 324313 168602 324379 168605
rect 248860 168600 252251 168602
rect 248860 168544 252190 168600
rect 252246 168544 252251 168600
rect 248860 168542 252251 168544
rect 321908 168600 324379 168602
rect 321908 168544 324318 168600
rect 324374 168544 324379 168600
rect 321908 168542 324379 168544
rect 252185 168539 252251 168542
rect 324313 168539 324379 168542
rect 307293 168466 307359 168469
rect 307293 168464 310132 168466
rect 307293 168408 307298 168464
rect 307354 168408 310132 168464
rect 307293 168406 310132 168408
rect 307293 168403 307359 168406
rect 214005 168330 214071 168333
rect 214005 168328 217212 168330
rect 214005 168272 214010 168328
rect 214066 168272 217212 168328
rect 214005 168270 217212 168272
rect 214005 168267 214071 168270
rect 265014 168194 265020 168196
rect 248860 168134 265020 168194
rect 265014 168132 265020 168134
rect 265084 168132 265090 168196
rect 307109 168058 307175 168061
rect 307109 168056 310132 168058
rect 307109 168000 307114 168056
rect 307170 168000 310132 168056
rect 307109 167998 310132 168000
rect 307109 167995 307175 167998
rect 324405 167786 324471 167789
rect 321908 167784 324471 167786
rect 321908 167728 324410 167784
rect 324466 167728 324471 167784
rect 321908 167726 324471 167728
rect 324405 167723 324471 167726
rect 213913 167650 213979 167653
rect 252461 167650 252527 167653
rect 213913 167648 217212 167650
rect 213913 167592 213918 167648
rect 213974 167592 217212 167648
rect 213913 167590 217212 167592
rect 248860 167648 252527 167650
rect 248860 167592 252466 167648
rect 252522 167592 252527 167648
rect 248860 167590 252527 167592
rect 213913 167587 213979 167590
rect 252461 167587 252527 167590
rect 306925 167650 306991 167653
rect 306925 167648 310132 167650
rect 306925 167592 306930 167648
rect 306986 167592 310132 167648
rect 306925 167590 310132 167592
rect 306925 167587 306991 167590
rect 252277 167242 252343 167245
rect 248860 167240 252343 167242
rect 248860 167184 252282 167240
rect 252338 167184 252343 167240
rect 248860 167182 252343 167184
rect 252277 167179 252343 167182
rect 307201 167242 307267 167245
rect 307201 167240 310132 167242
rect 307201 167184 307206 167240
rect 307262 167184 310132 167240
rect 307201 167182 310132 167184
rect 307201 167179 307267 167182
rect 324313 167106 324379 167109
rect 321908 167104 324379 167106
rect 321908 167048 324318 167104
rect 324374 167048 324379 167104
rect 321908 167046 324379 167048
rect 324313 167043 324379 167046
rect 213913 166970 213979 166973
rect 213913 166968 217212 166970
rect 213913 166912 213918 166968
rect 213974 166912 217212 166968
rect 213913 166910 217212 166912
rect 213913 166907 213979 166910
rect 306925 166834 306991 166837
rect 306925 166832 310132 166834
rect 306925 166776 306930 166832
rect 306986 166776 310132 166832
rect 306925 166774 310132 166776
rect 306925 166771 306991 166774
rect 252277 166698 252343 166701
rect 248860 166696 252343 166698
rect 248860 166640 252282 166696
rect 252338 166640 252343 166696
rect 248860 166638 252343 166640
rect 252277 166635 252343 166638
rect 214005 166426 214071 166429
rect 307661 166426 307727 166429
rect 214005 166424 217212 166426
rect 214005 166368 214010 166424
rect 214066 166368 217212 166424
rect 214005 166366 217212 166368
rect 307661 166424 310132 166426
rect 307661 166368 307666 166424
rect 307722 166368 310132 166424
rect 307661 166366 310132 166368
rect 214005 166363 214071 166366
rect 307661 166363 307727 166366
rect 251909 166290 251975 166293
rect 248860 166288 251975 166290
rect 248860 166232 251914 166288
rect 251970 166232 251975 166288
rect 248860 166230 251975 166232
rect 251909 166227 251975 166230
rect 307477 165882 307543 165885
rect 307477 165880 310132 165882
rect 307477 165824 307482 165880
rect 307538 165824 310132 165880
rect 307477 165822 310132 165824
rect 307477 165819 307543 165822
rect 213913 165746 213979 165749
rect 252277 165746 252343 165749
rect 213913 165744 217212 165746
rect 213913 165688 213918 165744
rect 213974 165688 217212 165744
rect 213913 165686 217212 165688
rect 248860 165744 252343 165746
rect 248860 165688 252282 165744
rect 252338 165688 252343 165744
rect 248860 165686 252343 165688
rect 321878 165746 321938 166260
rect 582557 165882 582623 165885
rect 583520 165882 584960 165972
rect 582557 165880 584960 165882
rect 582557 165824 582562 165880
rect 582618 165824 584960 165880
rect 582557 165822 584960 165824
rect 582557 165819 582623 165822
rect 334014 165746 334020 165748
rect 321878 165686 334020 165746
rect 213913 165683 213979 165686
rect 252277 165683 252343 165686
rect 334014 165684 334020 165686
rect 334084 165684 334090 165748
rect 583520 165732 584960 165822
rect 307569 165474 307635 165477
rect 324313 165474 324379 165477
rect 307569 165472 310132 165474
rect 307569 165416 307574 165472
rect 307630 165416 310132 165472
rect 307569 165414 310132 165416
rect 321908 165472 324379 165474
rect 321908 165416 324318 165472
rect 324374 165416 324379 165472
rect 321908 165414 324379 165416
rect 307569 165411 307635 165414
rect 324313 165411 324379 165414
rect 252461 165338 252527 165341
rect 248860 165336 252527 165338
rect 248860 165280 252466 165336
rect 252522 165280 252527 165336
rect 248860 165278 252527 165280
rect 252461 165275 252527 165278
rect 213913 165066 213979 165069
rect 307385 165066 307451 165069
rect 213913 165064 217212 165066
rect 213913 165008 213918 165064
rect 213974 165008 217212 165064
rect 213913 165006 217212 165008
rect 307385 165064 310132 165066
rect 307385 165008 307390 165064
rect 307446 165008 310132 165064
rect 307385 165006 310132 165008
rect 213913 165003 213979 165006
rect 307385 165003 307451 165006
rect 266302 164794 266308 164796
rect 248860 164734 266308 164794
rect 266302 164732 266308 164734
rect 266372 164732 266378 164796
rect 324405 164794 324471 164797
rect 321908 164792 324471 164794
rect 321908 164736 324410 164792
rect 324466 164736 324471 164792
rect 321908 164734 324471 164736
rect 324405 164731 324471 164734
rect 307661 164658 307727 164661
rect 307661 164656 310132 164658
rect 307661 164600 307666 164656
rect 307722 164600 310132 164656
rect 307661 164598 310132 164600
rect 307661 164595 307727 164598
rect 214005 164386 214071 164389
rect 251541 164386 251607 164389
rect 214005 164384 217212 164386
rect 214005 164328 214010 164384
rect 214066 164328 217212 164384
rect 214005 164326 217212 164328
rect 248860 164384 251607 164386
rect 248860 164328 251546 164384
rect 251602 164328 251607 164384
rect 248860 164326 251607 164328
rect 214005 164323 214071 164326
rect 251541 164323 251607 164326
rect 252829 164250 252895 164253
rect 256918 164250 256924 164252
rect 252829 164248 256924 164250
rect 252829 164192 252834 164248
rect 252890 164192 256924 164248
rect 252829 164190 256924 164192
rect 252829 164187 252895 164190
rect 256918 164188 256924 164190
rect 256988 164188 256994 164252
rect 307293 164250 307359 164253
rect 307293 164248 310132 164250
rect 307293 164192 307298 164248
rect 307354 164192 310132 164248
rect 307293 164190 310132 164192
rect 307293 164187 307359 164190
rect 252461 163978 252527 163981
rect 324313 163978 324379 163981
rect 248860 163976 252527 163978
rect 248860 163920 252466 163976
rect 252522 163920 252527 163976
rect 248860 163918 252527 163920
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 252461 163915 252527 163918
rect 324313 163915 324379 163918
rect 307569 163842 307635 163845
rect 307569 163840 310132 163842
rect 307569 163784 307574 163840
rect 307630 163784 310132 163840
rect 307569 163782 310132 163784
rect 307569 163779 307635 163782
rect 166390 163100 166396 163164
rect 166460 163162 166466 163164
rect 217182 163162 217242 163676
rect 263726 163434 263732 163436
rect 248860 163374 263732 163434
rect 263726 163372 263732 163374
rect 263796 163372 263802 163436
rect 307293 163434 307359 163437
rect 307293 163432 310132 163434
rect 307293 163376 307298 163432
rect 307354 163376 310132 163432
rect 307293 163374 310132 163376
rect 307293 163371 307359 163374
rect 324405 163162 324471 163165
rect 166460 163102 217242 163162
rect 321908 163160 324471 163162
rect 321908 163104 324410 163160
rect 324466 163104 324471 163160
rect 321908 163102 324471 163104
rect 166460 163100 166466 163102
rect 324405 163099 324471 163102
rect 213913 163026 213979 163029
rect 252093 163026 252159 163029
rect 213913 163024 217212 163026
rect 213913 162968 213918 163024
rect 213974 162968 217212 163024
rect 213913 162966 217212 162968
rect 248860 163024 252159 163026
rect 248860 162968 252098 163024
rect 252154 162968 252159 163024
rect 248860 162966 252159 162968
rect 213913 162963 213979 162966
rect 252093 162963 252159 162966
rect 307661 163026 307727 163029
rect 307661 163024 310132 163026
rect 307661 162968 307666 163024
rect 307722 162968 310132 163024
rect 307661 162966 310132 162968
rect 307661 162963 307727 162966
rect 305637 162890 305703 162893
rect 307569 162890 307635 162893
rect 305637 162888 307635 162890
rect 305637 162832 305642 162888
rect 305698 162832 307574 162888
rect 307630 162832 307635 162888
rect 305637 162830 307635 162832
rect 305637 162827 305703 162830
rect 307569 162827 307635 162830
rect 252461 162482 252527 162485
rect 248860 162480 252527 162482
rect 248860 162424 252466 162480
rect 252522 162424 252527 162480
rect 248860 162422 252527 162424
rect 252461 162419 252527 162422
rect 307477 162482 307543 162485
rect 307477 162480 310132 162482
rect 307477 162424 307482 162480
rect 307538 162424 310132 162480
rect 307477 162422 310132 162424
rect 307477 162419 307543 162422
rect 217182 161938 217242 162316
rect 252461 162074 252527 162077
rect 248860 162072 252527 162074
rect 248860 162016 252466 162072
rect 252522 162016 252527 162072
rect 248860 162014 252527 162016
rect 252461 162011 252527 162014
rect 307661 162074 307727 162077
rect 307661 162072 310132 162074
rect 307661 162016 307666 162072
rect 307722 162016 310132 162072
rect 307661 162014 310132 162016
rect 307661 162011 307727 162014
rect 200070 161878 217242 161938
rect 167678 161468 167684 161532
rect 167748 161530 167754 161532
rect 200070 161530 200130 161878
rect 214649 161802 214715 161805
rect 321878 161802 321938 162452
rect 214649 161800 217212 161802
rect 214649 161744 214654 161800
rect 214710 161744 217212 161800
rect 214649 161742 217212 161744
rect 321878 161742 325710 161802
rect 214649 161739 214715 161742
rect 307017 161666 307083 161669
rect 324313 161666 324379 161669
rect 307017 161664 310132 161666
rect 307017 161608 307022 161664
rect 307078 161608 310132 161664
rect 307017 161606 310132 161608
rect 321908 161664 324379 161666
rect 321908 161608 324318 161664
rect 324374 161608 324379 161664
rect 321908 161606 324379 161608
rect 307017 161603 307083 161606
rect 324313 161603 324379 161606
rect 252461 161530 252527 161533
rect 167748 161470 200130 161530
rect 248860 161528 252527 161530
rect 248860 161472 252466 161528
rect 252522 161472 252527 161528
rect 248860 161470 252527 161472
rect 325650 161530 325710 161742
rect 345054 161530 345060 161532
rect 325650 161470 345060 161530
rect 167748 161468 167754 161470
rect 252461 161467 252527 161470
rect 345054 161468 345060 161470
rect 345124 161468 345130 161532
rect 306741 161258 306807 161261
rect 306741 161256 310132 161258
rect 306741 161200 306746 161256
rect 306802 161200 310132 161256
rect 306741 161198 310132 161200
rect 306741 161195 306807 161198
rect 215017 161122 215083 161125
rect 252461 161122 252527 161125
rect 215017 161120 217212 161122
rect 215017 161064 215022 161120
rect 215078 161064 217212 161120
rect 215017 161062 217212 161064
rect 248860 161120 252527 161122
rect 248860 161064 252466 161120
rect 252522 161064 252527 161120
rect 248860 161062 252527 161064
rect 215017 161059 215083 161062
rect 252461 161059 252527 161062
rect 307477 160850 307543 160853
rect 307477 160848 310132 160850
rect 307477 160792 307482 160848
rect 307538 160792 310132 160848
rect 307477 160790 310132 160792
rect 307477 160787 307543 160790
rect 252737 160578 252803 160581
rect 248860 160576 252803 160578
rect 248860 160520 252742 160576
rect 252798 160520 252803 160576
rect 248860 160518 252803 160520
rect 252737 160515 252803 160518
rect 214925 160442 214991 160445
rect 307661 160442 307727 160445
rect 214925 160440 217212 160442
rect 214925 160384 214930 160440
rect 214986 160384 217212 160440
rect 214925 160382 217212 160384
rect 307661 160440 310132 160442
rect 307661 160384 307666 160440
rect 307722 160384 310132 160440
rect 307661 160382 310132 160384
rect 214925 160379 214991 160382
rect 307661 160379 307727 160382
rect 321878 160306 321938 160820
rect 321878 160246 325710 160306
rect 252461 160170 252527 160173
rect 324313 160170 324379 160173
rect 248860 160168 252527 160170
rect 248860 160112 252466 160168
rect 252522 160112 252527 160168
rect 248860 160110 252527 160112
rect 321908 160168 324379 160170
rect 321908 160112 324318 160168
rect 324374 160112 324379 160168
rect 321908 160110 324379 160112
rect 325650 160170 325710 160246
rect 335670 160170 335676 160172
rect 325650 160110 335676 160170
rect 252461 160107 252527 160110
rect 324313 160107 324379 160110
rect 335670 160108 335676 160110
rect 335740 160108 335746 160172
rect 307569 160034 307635 160037
rect 307569 160032 310132 160034
rect 307569 159976 307574 160032
rect 307630 159976 310132 160032
rect 307569 159974 310132 159976
rect 307569 159971 307635 159974
rect 213913 159762 213979 159765
rect 213913 159760 217212 159762
rect 213913 159704 213918 159760
rect 213974 159704 217212 159760
rect 213913 159702 217212 159704
rect 213913 159699 213979 159702
rect 252461 159626 252527 159629
rect 248860 159624 252527 159626
rect 248860 159568 252466 159624
rect 252522 159568 252527 159624
rect 248860 159566 252527 159568
rect 252461 159563 252527 159566
rect 307661 159626 307727 159629
rect 307661 159624 310132 159626
rect 307661 159568 307666 159624
rect 307722 159568 310132 159624
rect 307661 159566 310132 159568
rect 307661 159563 307727 159566
rect 324313 159354 324379 159357
rect 321908 159352 324379 159354
rect 321908 159296 324318 159352
rect 324374 159296 324379 159352
rect 321908 159294 324379 159296
rect 324313 159291 324379 159294
rect 251909 159218 251975 159221
rect 248860 159216 251975 159218
rect 248860 159160 251914 159216
rect 251970 159160 251975 159216
rect 248860 159158 251975 159160
rect 251909 159155 251975 159158
rect 214005 159082 214071 159085
rect 307201 159082 307267 159085
rect 214005 159080 217212 159082
rect 214005 159024 214010 159080
rect 214066 159024 217212 159080
rect 214005 159022 217212 159024
rect 307201 159080 310132 159082
rect 307201 159024 307206 159080
rect 307262 159024 310132 159080
rect 307201 159022 310132 159024
rect 214005 159019 214071 159022
rect 307201 159019 307267 159022
rect 251449 158810 251515 158813
rect 248860 158808 251515 158810
rect 248860 158752 251454 158808
rect 251510 158752 251515 158808
rect 248860 158750 251515 158752
rect 251449 158747 251515 158750
rect 306925 158674 306991 158677
rect 306925 158672 310132 158674
rect 306925 158616 306930 158672
rect 306986 158616 310132 158672
rect 306925 158614 310132 158616
rect 306925 158611 306991 158614
rect 324313 158538 324379 158541
rect 321908 158536 324379 158538
rect 321908 158480 324318 158536
rect 324374 158480 324379 158536
rect 321908 158478 324379 158480
rect 324313 158475 324379 158478
rect 217182 157858 217242 158372
rect 252461 158266 252527 158269
rect 248860 158264 252527 158266
rect 248860 158208 252466 158264
rect 252522 158208 252527 158264
rect 248860 158206 252527 158208
rect 252461 158203 252527 158206
rect 307661 158266 307727 158269
rect 307661 158264 310132 158266
rect 307661 158208 307666 158264
rect 307722 158208 310132 158264
rect 307661 158206 310132 158208
rect 307661 158203 307727 158206
rect 262254 157858 262260 157860
rect 200070 157798 217242 157858
rect 248860 157798 262260 157858
rect 167494 157388 167500 157452
rect 167564 157450 167570 157452
rect 200070 157450 200130 157798
rect 262254 157796 262260 157798
rect 262324 157796 262330 157860
rect 307293 157858 307359 157861
rect 324405 157858 324471 157861
rect 307293 157856 310132 157858
rect 307293 157800 307298 157856
rect 307354 157800 310132 157856
rect 307293 157798 310132 157800
rect 321908 157856 324471 157858
rect 321908 157800 324410 157856
rect 324466 157800 324471 157856
rect 321908 157798 324471 157800
rect 307293 157795 307359 157798
rect 324405 157795 324471 157798
rect 213913 157722 213979 157725
rect 213913 157720 217212 157722
rect 213913 157664 213918 157720
rect 213974 157664 217212 157720
rect 213913 157662 217212 157664
rect 213913 157659 213979 157662
rect 167564 157390 200130 157450
rect 307661 157450 307727 157453
rect 307661 157448 310132 157450
rect 307661 157392 307666 157448
rect 307722 157392 310132 157448
rect 307661 157390 310132 157392
rect 167564 157388 167570 157390
rect 307661 157387 307727 157390
rect 252461 157314 252527 157317
rect 248860 157312 252527 157314
rect 248860 157256 252466 157312
rect 252522 157256 252527 157312
rect 248860 157254 252527 157256
rect 252461 157251 252527 157254
rect 213913 157178 213979 157181
rect 213913 157176 217212 157178
rect 213913 157120 213918 157176
rect 213974 157120 217212 157176
rect 213913 157118 217212 157120
rect 213913 157115 213979 157118
rect 306741 157042 306807 157045
rect 324313 157042 324379 157045
rect 306741 157040 310132 157042
rect 306741 156984 306746 157040
rect 306802 156984 310132 157040
rect 306741 156982 310132 156984
rect 321908 157040 324379 157042
rect 321908 156984 324318 157040
rect 324374 156984 324379 157040
rect 321908 156982 324379 156984
rect 306741 156979 306807 156982
rect 324313 156979 324379 156982
rect 251541 156906 251607 156909
rect 248860 156904 251607 156906
rect 248860 156848 251546 156904
rect 251602 156848 251607 156904
rect 248860 156846 251607 156848
rect 251541 156843 251607 156846
rect 307477 156634 307543 156637
rect 307477 156632 310132 156634
rect 307477 156576 307482 156632
rect 307538 156576 310132 156632
rect 307477 156574 310132 156576
rect 307477 156571 307543 156574
rect 214005 156498 214071 156501
rect 214005 156496 217212 156498
rect 214005 156440 214010 156496
rect 214066 156440 217212 156496
rect 214005 156438 217212 156440
rect 214005 156435 214071 156438
rect 251357 156362 251423 156365
rect 324405 156362 324471 156365
rect 248860 156360 251423 156362
rect 248860 156304 251362 156360
rect 251418 156304 251423 156360
rect 248860 156302 251423 156304
rect 321908 156360 324471 156362
rect 321908 156304 324410 156360
rect 324466 156304 324471 156360
rect 321908 156302 324471 156304
rect 251357 156299 251423 156302
rect 324405 156299 324471 156302
rect 307385 156226 307451 156229
rect 307385 156224 310132 156226
rect 307385 156168 307390 156224
rect 307446 156168 310132 156224
rect 307385 156166 310132 156168
rect 307385 156163 307451 156166
rect 252461 155954 252527 155957
rect 248860 155952 252527 155954
rect 248860 155896 252466 155952
rect 252522 155896 252527 155952
rect 248860 155894 252527 155896
rect 252461 155891 252527 155894
rect 213913 155818 213979 155821
rect 213913 155816 217212 155818
rect 213913 155760 213918 155816
rect 213974 155760 217212 155816
rect 213913 155758 217212 155760
rect 213913 155755 213979 155758
rect 307477 155682 307543 155685
rect 307477 155680 310132 155682
rect 307477 155624 307482 155680
rect 307538 155624 310132 155680
rect 307477 155622 310132 155624
rect 307477 155619 307543 155622
rect 324589 155546 324655 155549
rect 321908 155544 324655 155546
rect 321908 155488 324594 155544
rect 324650 155488 324655 155544
rect 321908 155486 324655 155488
rect 324589 155483 324655 155486
rect 252502 155410 252508 155412
rect 248860 155350 252508 155410
rect 252502 155348 252508 155350
rect 252572 155348 252578 155412
rect 307569 155274 307635 155277
rect 307569 155272 310132 155274
rect 307569 155216 307574 155272
rect 307630 155216 310132 155272
rect 307569 155214 310132 155216
rect 307569 155211 307635 155214
rect 166206 154532 166212 154596
rect 166276 154594 166282 154596
rect 217182 154594 217242 155108
rect 252369 155002 252435 155005
rect 248860 155000 252435 155002
rect 248860 154944 252374 155000
rect 252430 154944 252435 155000
rect 248860 154942 252435 154944
rect 252369 154939 252435 154942
rect 307661 154866 307727 154869
rect 307661 154864 310132 154866
rect 307661 154808 307666 154864
rect 307722 154808 310132 154864
rect 307661 154806 310132 154808
rect 307661 154803 307727 154806
rect 324313 154730 324379 154733
rect 321908 154728 324379 154730
rect 321908 154672 324318 154728
rect 324374 154672 324379 154728
rect 321908 154670 324379 154672
rect 324313 154667 324379 154670
rect 166276 154534 217242 154594
rect 166276 154532 166282 154534
rect 214005 154458 214071 154461
rect 252461 154458 252527 154461
rect 214005 154456 217212 154458
rect 214005 154400 214010 154456
rect 214066 154400 217212 154456
rect 214005 154398 217212 154400
rect 248860 154456 252527 154458
rect 248860 154400 252466 154456
rect 252522 154400 252527 154456
rect 248860 154398 252527 154400
rect 214005 154395 214071 154398
rect 252461 154395 252527 154398
rect 307477 154458 307543 154461
rect 307477 154456 310132 154458
rect 307477 154400 307482 154456
rect 307538 154400 310132 154456
rect 307477 154398 310132 154400
rect 307477 154395 307543 154398
rect 251541 154050 251607 154053
rect 248860 154048 251607 154050
rect 248860 153992 251546 154048
rect 251602 153992 251607 154048
rect 248860 153990 251607 153992
rect 251541 153987 251607 153990
rect 307661 154050 307727 154053
rect 324313 154050 324379 154053
rect 307661 154048 310132 154050
rect 307661 153992 307666 154048
rect 307722 153992 310132 154048
rect 307661 153990 310132 153992
rect 321908 154048 324379 154050
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 307661 153987 307727 153990
rect 324313 153987 324379 153990
rect 213913 153778 213979 153781
rect 213913 153776 217212 153778
rect 213913 153720 213918 153776
rect 213974 153720 217212 153776
rect 213913 153718 217212 153720
rect 213913 153715 213979 153718
rect 307569 153642 307635 153645
rect 307569 153640 310132 153642
rect 307569 153584 307574 153640
rect 307630 153584 310132 153640
rect 307569 153582 310132 153584
rect 307569 153579 307635 153582
rect 252001 153506 252067 153509
rect 248860 153504 252067 153506
rect 248860 153448 252006 153504
rect 252062 153448 252067 153504
rect 248860 153446 252067 153448
rect 252001 153443 252067 153446
rect 306649 153234 306715 153237
rect 324405 153234 324471 153237
rect 306649 153232 310132 153234
rect 306649 153176 306654 153232
rect 306710 153176 310132 153232
rect 306649 153174 310132 153176
rect 321908 153232 324471 153234
rect 321908 153176 324410 153232
rect 324466 153176 324471 153232
rect 321908 153174 324471 153176
rect 306649 153171 306715 153174
rect 324405 153171 324471 153174
rect 214005 153098 214071 153101
rect 252461 153098 252527 153101
rect 214005 153096 217212 153098
rect 214005 153040 214010 153096
rect 214066 153040 217212 153096
rect 214005 153038 217212 153040
rect 248860 153096 252527 153098
rect 248860 153040 252466 153096
rect 252522 153040 252527 153096
rect 248860 153038 252527 153040
rect 214005 153035 214071 153038
rect 252461 153035 252527 153038
rect 252277 152690 252343 152693
rect 248860 152688 252343 152690
rect 248860 152632 252282 152688
rect 252338 152632 252343 152688
rect 248860 152630 252343 152632
rect 252277 152627 252343 152630
rect 307477 152690 307543 152693
rect 582373 152690 582439 152693
rect 583520 152690 584960 152780
rect 307477 152688 310132 152690
rect 307477 152632 307482 152688
rect 307538 152632 310132 152688
rect 307477 152630 310132 152632
rect 582373 152688 584960 152690
rect 582373 152632 582378 152688
rect 582434 152632 584960 152688
rect 582373 152630 584960 152632
rect 307477 152627 307543 152630
rect 582373 152627 582439 152630
rect 213913 152554 213979 152557
rect 213913 152552 217212 152554
rect 213913 152496 213918 152552
rect 213974 152496 217212 152552
rect 583520 152540 584960 152630
rect 213913 152494 217212 152496
rect 213913 152491 213979 152494
rect 324313 152418 324379 152421
rect 321908 152416 324379 152418
rect 321908 152360 324318 152416
rect 324374 152360 324379 152416
rect 321908 152358 324379 152360
rect 324313 152355 324379 152358
rect 306557 152282 306623 152285
rect 306557 152280 310132 152282
rect 306557 152224 306562 152280
rect 306618 152224 310132 152280
rect 306557 152222 310132 152224
rect 306557 152219 306623 152222
rect 251725 152146 251791 152149
rect 248860 152144 251791 152146
rect 248860 152088 251730 152144
rect 251786 152088 251791 152144
rect 248860 152086 251791 152088
rect 251725 152083 251791 152086
rect 214649 151874 214715 151877
rect 307661 151874 307727 151877
rect 214649 151872 217212 151874
rect 214649 151816 214654 151872
rect 214710 151816 217212 151872
rect 214649 151814 217212 151816
rect 307661 151872 310132 151874
rect 307661 151816 307666 151872
rect 307722 151816 310132 151872
rect 307661 151814 310132 151816
rect 214649 151811 214715 151814
rect 307661 151811 307727 151814
rect 252461 151738 252527 151741
rect 324313 151738 324379 151741
rect 248860 151736 252527 151738
rect 248860 151680 252466 151736
rect 252522 151680 252527 151736
rect 248860 151678 252527 151680
rect 321908 151736 324379 151738
rect 321908 151680 324318 151736
rect 324374 151680 324379 151736
rect 321908 151678 324379 151680
rect 252461 151675 252527 151678
rect 324313 151675 324379 151678
rect 307477 151466 307543 151469
rect 307477 151464 310132 151466
rect 307477 151408 307482 151464
rect 307538 151408 310132 151464
rect 307477 151406 310132 151408
rect 307477 151403 307543 151406
rect 214097 151194 214163 151197
rect 251265 151194 251331 151197
rect 214097 151192 217212 151194
rect 214097 151136 214102 151192
rect 214158 151136 217212 151192
rect 214097 151134 217212 151136
rect 248860 151192 251331 151194
rect 248860 151136 251270 151192
rect 251326 151136 251331 151192
rect 248860 151134 251331 151136
rect 214097 151131 214163 151134
rect 251265 151131 251331 151134
rect 307661 151058 307727 151061
rect 307661 151056 310132 151058
rect 307661 151000 307666 151056
rect 307722 151000 310132 151056
rect 307661 150998 310132 151000
rect 307661 150995 307727 150998
rect 324405 150922 324471 150925
rect 321908 150920 324471 150922
rect 321908 150864 324410 150920
rect 324466 150864 324471 150920
rect 321908 150862 324471 150864
rect 324405 150859 324471 150862
rect 252369 150786 252435 150789
rect 248860 150784 252435 150786
rect 248860 150728 252374 150784
rect 252430 150728 252435 150784
rect 248860 150726 252435 150728
rect 252369 150723 252435 150726
rect 307385 150650 307451 150653
rect 307385 150648 310132 150650
rect 307385 150592 307390 150648
rect 307446 150592 310132 150648
rect 307385 150590 310132 150592
rect 307385 150587 307451 150590
rect 213913 150514 213979 150517
rect 213913 150512 217212 150514
rect 213913 150456 213918 150512
rect 213974 150456 217212 150512
rect 213913 150454 217212 150456
rect 213913 150451 213979 150454
rect 322054 150378 322060 150380
rect 321878 150318 322060 150378
rect 252461 150242 252527 150245
rect 248860 150240 252527 150242
rect 248860 150184 252466 150240
rect 252522 150184 252527 150240
rect 248860 150182 252527 150184
rect 252461 150179 252527 150182
rect 306925 150242 306991 150245
rect 306925 150240 310132 150242
rect 306925 150184 306930 150240
rect 306986 150184 310132 150240
rect 306925 150182 310132 150184
rect 306925 150179 306991 150182
rect 321878 150076 321938 150318
rect 322054 150316 322060 150318
rect 322124 150316 322130 150380
rect 214557 149834 214623 149837
rect 249885 149834 249951 149837
rect 214557 149832 217212 149834
rect 214557 149776 214562 149832
rect 214618 149776 217212 149832
rect 214557 149774 217212 149776
rect 248860 149832 249951 149834
rect 248860 149776 249890 149832
rect 249946 149776 249951 149832
rect 248860 149774 249951 149776
rect 214557 149771 214623 149774
rect 249885 149771 249951 149774
rect 307477 149834 307543 149837
rect 307477 149832 310132 149834
rect 307477 149776 307482 149832
rect 307538 149776 310132 149832
rect 307477 149774 310132 149776
rect 307477 149771 307543 149774
rect 324313 149426 324379 149429
rect 321908 149424 324379 149426
rect 321908 149368 324318 149424
rect 324374 149368 324379 149424
rect 321908 149366 324379 149368
rect 324313 149363 324379 149366
rect 251725 149290 251791 149293
rect 248860 149288 251791 149290
rect 248860 149232 251730 149288
rect 251786 149232 251791 149288
rect 248860 149230 251791 149232
rect 251725 149227 251791 149230
rect 307293 149290 307359 149293
rect 307293 149288 310132 149290
rect 307293 149232 307298 149288
rect 307354 149232 310132 149288
rect 307293 149230 310132 149232
rect 307293 149227 307359 149230
rect 214005 149154 214071 149157
rect 214005 149152 217212 149154
rect 214005 149096 214010 149152
rect 214066 149096 217212 149152
rect 214005 149094 217212 149096
rect 214005 149091 214071 149094
rect 252461 148882 252527 148885
rect 248860 148880 252527 148882
rect 248860 148824 252466 148880
rect 252522 148824 252527 148880
rect 248860 148822 252527 148824
rect 252461 148819 252527 148822
rect 307661 148882 307727 148885
rect 307661 148880 310132 148882
rect 307661 148824 307666 148880
rect 307722 148824 310132 148880
rect 307661 148822 310132 148824
rect 307661 148819 307727 148822
rect 324313 148610 324379 148613
rect 321908 148608 324379 148610
rect 321908 148552 324318 148608
rect 324374 148552 324379 148608
rect 321908 148550 324379 148552
rect 324313 148547 324379 148550
rect 213913 148474 213979 148477
rect 307477 148474 307543 148477
rect 213913 148472 217212 148474
rect 213913 148416 213918 148472
rect 213974 148416 217212 148472
rect 213913 148414 217212 148416
rect 307477 148472 310132 148474
rect 307477 148416 307482 148472
rect 307538 148416 310132 148472
rect 307477 148414 310132 148416
rect 213913 148411 213979 148414
rect 307477 148411 307543 148414
rect 251541 148338 251607 148341
rect 248860 148336 251607 148338
rect 248860 148280 251546 148336
rect 251602 148280 251607 148336
rect 248860 148278 251607 148280
rect 251541 148275 251607 148278
rect 321645 148338 321711 148341
rect 321645 148336 321754 148338
rect 321645 148280 321650 148336
rect 321706 148280 321754 148336
rect 321645 148275 321754 148280
rect 307109 148066 307175 148069
rect 307109 148064 310132 148066
rect 307109 148008 307114 148064
rect 307170 148008 310132 148064
rect 307109 148006 310132 148008
rect 307109 148003 307175 148006
rect 213913 147930 213979 147933
rect 255446 147930 255452 147932
rect 213913 147928 217212 147930
rect 213913 147872 213918 147928
rect 213974 147872 217212 147928
rect 213913 147870 217212 147872
rect 248860 147870 255452 147930
rect 213913 147867 213979 147870
rect 255446 147868 255452 147870
rect 255516 147868 255522 147932
rect 321694 147764 321754 148275
rect 307293 147658 307359 147661
rect 307293 147656 310132 147658
rect 307293 147600 307298 147656
rect 307354 147600 310132 147656
rect 307293 147598 310132 147600
rect 307293 147595 307359 147598
rect 252461 147522 252527 147525
rect 248860 147520 252527 147522
rect 248860 147464 252466 147520
rect 252522 147464 252527 147520
rect 248860 147462 252527 147464
rect 252461 147459 252527 147462
rect 213913 147250 213979 147253
rect 306741 147250 306807 147253
rect 213913 147248 217212 147250
rect 213913 147192 213918 147248
rect 213974 147192 217212 147248
rect 213913 147190 217212 147192
rect 306741 147248 310132 147250
rect 306741 147192 306746 147248
rect 306802 147192 310132 147248
rect 306741 147190 310132 147192
rect 213913 147187 213979 147190
rect 306741 147187 306807 147190
rect 324313 147114 324379 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 324313 147051 324379 147054
rect 251265 146978 251331 146981
rect 248860 146976 251331 146978
rect 248860 146920 251270 146976
rect 251326 146920 251331 146976
rect 248860 146918 251331 146920
rect 251265 146915 251331 146918
rect 307661 146842 307727 146845
rect 307661 146840 310132 146842
rect 307661 146784 307666 146840
rect 307722 146784 310132 146840
rect 307661 146782 310132 146784
rect 307661 146779 307727 146782
rect 214557 146570 214623 146573
rect 251357 146570 251423 146573
rect 214557 146568 217212 146570
rect 214557 146512 214562 146568
rect 214618 146512 217212 146568
rect 214557 146510 217212 146512
rect 248860 146568 251423 146570
rect 248860 146512 251362 146568
rect 251418 146512 251423 146568
rect 248860 146510 251423 146512
rect 214557 146507 214623 146510
rect 251357 146507 251423 146510
rect 307569 146434 307635 146437
rect 307569 146432 310132 146434
rect 307569 146376 307574 146432
rect 307630 146376 310132 146432
rect 307569 146374 310132 146376
rect 307569 146371 307635 146374
rect 251725 146298 251791 146301
rect 257838 146298 257844 146300
rect 251725 146296 257844 146298
rect 251725 146240 251730 146296
rect 251786 146240 257844 146296
rect 251725 146238 257844 146240
rect 251725 146235 251791 146238
rect 257838 146236 257844 146238
rect 257908 146236 257914 146300
rect 323669 146298 323735 146301
rect 321908 146296 323735 146298
rect 321908 146240 323674 146296
rect 323730 146240 323735 146296
rect 321908 146238 323735 146240
rect 323669 146235 323735 146238
rect 252461 146026 252527 146029
rect 248860 146024 252527 146026
rect 248860 145968 252466 146024
rect 252522 145968 252527 146024
rect 248860 145966 252527 145968
rect 252461 145963 252527 145966
rect 213913 145890 213979 145893
rect 307477 145890 307543 145893
rect 213913 145888 217212 145890
rect 213913 145832 213918 145888
rect 213974 145832 217212 145888
rect 213913 145830 217212 145832
rect 307477 145888 310132 145890
rect 307477 145832 307482 145888
rect 307538 145832 310132 145888
rect 307477 145830 310132 145832
rect 213913 145827 213979 145830
rect 307477 145827 307543 145830
rect 252369 145618 252435 145621
rect 248860 145616 252435 145618
rect 248860 145560 252374 145616
rect 252430 145560 252435 145616
rect 248860 145558 252435 145560
rect 252369 145555 252435 145558
rect 307201 145482 307267 145485
rect 325785 145482 325851 145485
rect 307201 145480 310132 145482
rect 307201 145424 307206 145480
rect 307262 145424 310132 145480
rect 307201 145422 310132 145424
rect 321908 145480 325851 145482
rect 321908 145424 325790 145480
rect 325846 145424 325851 145480
rect 321908 145422 325851 145424
rect 307201 145419 307267 145422
rect 325785 145419 325851 145422
rect 214465 145210 214531 145213
rect 214465 145208 217212 145210
rect 214465 145152 214470 145208
rect 214526 145152 217212 145208
rect 214465 145150 217212 145152
rect 214465 145147 214531 145150
rect 252093 145074 252159 145077
rect 248860 145072 252159 145074
rect 248860 145016 252098 145072
rect 252154 145016 252159 145072
rect 248860 145014 252159 145016
rect 252093 145011 252159 145014
rect 307661 145074 307727 145077
rect 307661 145072 310132 145074
rect 307661 145016 307666 145072
rect 307722 145016 310132 145072
rect 307661 145014 310132 145016
rect 307661 145011 307727 145014
rect 324313 144802 324379 144805
rect 321908 144800 324379 144802
rect 321908 144744 324318 144800
rect 324374 144744 324379 144800
rect 321908 144742 324379 144744
rect 324313 144739 324379 144742
rect 252461 144666 252527 144669
rect 248860 144664 252527 144666
rect 248860 144608 252466 144664
rect 252522 144608 252527 144664
rect 248860 144606 252527 144608
rect 252461 144603 252527 144606
rect 306925 144666 306991 144669
rect 306925 144664 310132 144666
rect 306925 144608 306930 144664
rect 306986 144608 310132 144664
rect 306925 144606 310132 144608
rect 306925 144603 306991 144606
rect 213913 144530 213979 144533
rect 213913 144528 217212 144530
rect 213913 144472 213918 144528
rect 213974 144472 217212 144528
rect 213913 144470 217212 144472
rect 213913 144467 213979 144470
rect 306557 144258 306623 144261
rect 306557 144256 310132 144258
rect 306557 144200 306562 144256
rect 306618 144200 310132 144256
rect 306557 144198 310132 144200
rect 306557 144195 306623 144198
rect 251541 144122 251607 144125
rect 248860 144120 251607 144122
rect 248860 144064 251546 144120
rect 251602 144064 251607 144120
rect 248860 144062 251607 144064
rect 251541 144059 251607 144062
rect 307477 143850 307543 143853
rect 200070 143790 217212 143850
rect 307477 143848 310132 143850
rect 307477 143792 307482 143848
rect 307538 143792 310132 143848
rect 307477 143790 310132 143792
rect 167494 143652 167500 143716
rect 167564 143714 167570 143716
rect 200070 143714 200130 143790
rect 307477 143787 307543 143790
rect 252093 143714 252159 143717
rect 167564 143654 200130 143714
rect 248860 143712 252159 143714
rect 248860 143656 252098 143712
rect 252154 143656 252159 143712
rect 248860 143654 252159 143656
rect 167564 143652 167570 143654
rect 252093 143651 252159 143654
rect 321878 143578 321938 143956
rect 329782 143578 329788 143580
rect 321878 143518 329788 143578
rect 329782 143516 329788 143518
rect 329852 143516 329858 143580
rect 307661 143442 307727 143445
rect 307661 143440 310132 143442
rect 307661 143384 307666 143440
rect 307722 143384 310132 143440
rect 307661 143382 310132 143384
rect 307661 143379 307727 143382
rect 213913 143306 213979 143309
rect 213913 143304 217212 143306
rect 213913 143248 213918 143304
rect 213974 143248 217212 143304
rect 213913 143246 217212 143248
rect 213913 143243 213979 143246
rect 251725 143170 251791 143173
rect 324313 143170 324379 143173
rect 248860 143168 251791 143170
rect 248860 143112 251730 143168
rect 251786 143112 251791 143168
rect 248860 143110 251791 143112
rect 321908 143168 324379 143170
rect 321908 143112 324318 143168
rect 324374 143112 324379 143168
rect 321908 143110 324379 143112
rect 251725 143107 251791 143110
rect 324313 143107 324379 143110
rect 306741 143034 306807 143037
rect 306741 143032 310132 143034
rect 306741 142976 306746 143032
rect 306802 142976 310132 143032
rect 306741 142974 310132 142976
rect 306741 142971 306807 142974
rect 260966 142762 260972 142764
rect 248860 142702 260972 142762
rect 260966 142700 260972 142702
rect 261036 142700 261042 142764
rect 214925 142626 214991 142629
rect 214925 142624 217212 142626
rect 214925 142568 214930 142624
rect 214986 142568 217212 142624
rect 214925 142566 217212 142568
rect 214925 142563 214991 142566
rect 307293 142490 307359 142493
rect 307293 142488 310132 142490
rect 307293 142432 307298 142488
rect 307354 142432 310132 142488
rect 307293 142430 310132 142432
rect 307293 142427 307359 142430
rect 263542 142218 263548 142220
rect 248860 142158 263548 142218
rect 263542 142156 263548 142158
rect 263612 142156 263618 142220
rect 321878 142218 321938 142460
rect 328678 142218 328684 142220
rect 321878 142158 328684 142218
rect 328678 142156 328684 142158
rect 328748 142156 328754 142220
rect 307569 142082 307635 142085
rect 327165 142082 327231 142085
rect 328494 142082 328500 142084
rect 307569 142080 310132 142082
rect 307569 142024 307574 142080
rect 307630 142024 310132 142080
rect 307569 142022 310132 142024
rect 321878 142080 328500 142082
rect 321878 142024 327170 142080
rect 327226 142024 328500 142080
rect 321878 142022 328500 142024
rect 307569 142019 307635 142022
rect 213913 141946 213979 141949
rect 213913 141944 217212 141946
rect 213913 141888 213918 141944
rect 213974 141888 217212 141944
rect 213913 141886 217212 141888
rect 213913 141883 213979 141886
rect 252461 141810 252527 141813
rect 248860 141808 252527 141810
rect 248860 141752 252466 141808
rect 252522 141752 252527 141808
rect 248860 141750 252527 141752
rect 252461 141747 252527 141750
rect 307477 141674 307543 141677
rect 307477 141672 310132 141674
rect 307477 141616 307482 141672
rect 307538 141616 310132 141672
rect 321878 141644 321938 142022
rect 327165 142019 327231 142022
rect 328494 142020 328500 142022
rect 328564 142020 328570 142084
rect 307477 141614 310132 141616
rect 307477 141611 307543 141614
rect 252369 141538 252435 141541
rect 261334 141538 261340 141540
rect 252369 141536 261340 141538
rect 252369 141480 252374 141536
rect 252430 141480 261340 141536
rect 252369 141478 261340 141480
rect 252369 141475 252435 141478
rect 261334 141476 261340 141478
rect 261404 141476 261410 141540
rect 252829 141402 252895 141405
rect 269941 141402 270007 141405
rect 248860 141342 252754 141402
rect 213177 141266 213243 141269
rect 252694 141266 252754 141342
rect 252829 141400 270007 141402
rect 252829 141344 252834 141400
rect 252890 141344 269946 141400
rect 270002 141344 270007 141400
rect 252829 141342 270007 141344
rect 252829 141339 252895 141342
rect 269941 141339 270007 141342
rect 259678 141266 259684 141268
rect 213177 141264 217212 141266
rect 213177 141208 213182 141264
rect 213238 141208 217212 141264
rect 213177 141206 217212 141208
rect 252694 141206 259684 141266
rect 213177 141203 213243 141206
rect 259678 141204 259684 141206
rect 259748 141204 259754 141268
rect 307017 141266 307083 141269
rect 307017 141264 310132 141266
rect 307017 141208 307022 141264
rect 307078 141208 310132 141264
rect 307017 141206 310132 141208
rect 307017 141203 307083 141206
rect 251766 141068 251772 141132
rect 251836 141130 251842 141132
rect 252829 141130 252895 141133
rect 251836 141128 252895 141130
rect 251836 141072 252834 141128
rect 252890 141072 252895 141128
rect 251836 141070 252895 141072
rect 251836 141068 251842 141070
rect 252829 141067 252895 141070
rect 251173 140858 251239 140861
rect 248860 140856 251239 140858
rect 248860 140800 251178 140856
rect 251234 140800 251239 140856
rect 248860 140798 251239 140800
rect 251173 140795 251239 140798
rect 307661 140858 307727 140861
rect 336958 140858 336964 140860
rect 307661 140856 310132 140858
rect 307661 140800 307666 140856
rect 307722 140800 310132 140856
rect 307661 140798 310132 140800
rect 321908 140798 336964 140858
rect 307661 140795 307727 140798
rect 336958 140796 336964 140798
rect 337028 140796 337034 140860
rect 214005 140586 214071 140589
rect 214005 140584 217212 140586
rect 214005 140528 214010 140584
rect 214066 140528 217212 140584
rect 214005 140526 217212 140528
rect 214005 140523 214071 140526
rect 251173 140450 251239 140453
rect 248860 140448 251239 140450
rect 248860 140392 251178 140448
rect 251234 140392 251239 140448
rect 248860 140390 251239 140392
rect 251173 140387 251239 140390
rect 308262 140390 310132 140450
rect 253197 140042 253263 140045
rect 306966 140042 306972 140044
rect 253197 140040 306972 140042
rect 253197 139984 253202 140040
rect 253258 139984 306972 140040
rect 253197 139982 306972 139984
rect 253197 139979 253263 139982
rect 306966 139980 306972 139982
rect 307036 139980 307042 140044
rect 213913 139906 213979 139909
rect 255262 139906 255268 139908
rect 213913 139904 217212 139906
rect 213913 139848 213918 139904
rect 213974 139848 217212 139904
rect 213913 139846 217212 139848
rect 248860 139846 255268 139906
rect 213913 139843 213979 139846
rect 255262 139844 255268 139846
rect 255332 139844 255338 139908
rect 261334 139708 261340 139772
rect 261404 139770 261410 139772
rect 308262 139770 308322 140390
rect 308673 140042 308739 140045
rect 308673 140040 310132 140042
rect 308673 139984 308678 140040
rect 308734 139984 310132 140040
rect 308673 139982 310132 139984
rect 308673 139979 308739 139982
rect 261404 139710 308322 139770
rect 261404 139708 261410 139710
rect 307661 139634 307727 139637
rect 307661 139632 310132 139634
rect 307661 139576 307666 139632
rect 307722 139576 310132 139632
rect 307661 139574 310132 139576
rect 307661 139571 307727 139574
rect 249793 139498 249859 139501
rect 248860 139496 249859 139498
rect 248860 139440 249798 139496
rect 249854 139440 249859 139496
rect 248860 139438 249859 139440
rect 249793 139435 249859 139438
rect 305494 139436 305500 139500
rect 305564 139498 305570 139500
rect 308673 139498 308739 139501
rect 305564 139496 308739 139498
rect 305564 139440 308678 139496
rect 308734 139440 308739 139496
rect 305564 139438 308739 139440
rect 321878 139498 321938 140148
rect 346342 139498 346348 139500
rect 321878 139438 346348 139498
rect 305564 139436 305570 139438
rect 308673 139435 308739 139438
rect 346342 139436 346348 139438
rect 346412 139436 346418 139500
rect 327022 139362 327028 139364
rect 321908 139302 327028 139362
rect 327022 139300 327028 139302
rect 327092 139300 327098 139364
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 214005 139226 214071 139229
rect 214005 139224 217212 139226
rect 214005 139168 214010 139224
rect 214066 139168 217212 139224
rect 583520 139212 584960 139302
rect 214005 139166 217212 139168
rect 214005 139163 214071 139166
rect 307477 139090 307543 139093
rect 307477 139088 310132 139090
rect 307477 139032 307482 139088
rect 307538 139032 310132 139088
rect 307477 139030 310132 139032
rect 307477 139027 307543 139030
rect 259494 138954 259500 138956
rect 248860 138894 259500 138954
rect 259494 138892 259500 138894
rect 259564 138892 259570 138956
rect 213913 138682 213979 138685
rect 307569 138682 307635 138685
rect 213913 138680 217212 138682
rect 213913 138624 213918 138680
rect 213974 138624 217212 138680
rect 213913 138622 217212 138624
rect 307569 138680 310132 138682
rect 307569 138624 307574 138680
rect 307630 138624 310132 138680
rect 307569 138622 310132 138624
rect 213913 138619 213979 138622
rect 307569 138619 307635 138622
rect 252461 138546 252527 138549
rect 324313 138546 324379 138549
rect 248860 138544 252527 138546
rect 248860 138488 252466 138544
rect 252522 138488 252527 138544
rect 248860 138486 252527 138488
rect 321908 138544 324379 138546
rect 321908 138488 324318 138544
rect 324374 138488 324379 138544
rect 321908 138486 324379 138488
rect 252461 138483 252527 138486
rect 324313 138483 324379 138486
rect 307661 138274 307727 138277
rect 307661 138272 310132 138274
rect 307661 138216 307666 138272
rect 307722 138216 310132 138272
rect 307661 138214 310132 138216
rect 307661 138211 307727 138214
rect 214097 138002 214163 138005
rect 250805 138002 250871 138005
rect 214097 138000 217212 138002
rect 214097 137944 214102 138000
rect 214158 137944 217212 138000
rect 214097 137942 217212 137944
rect 248860 138000 250871 138002
rect 248860 137944 250810 138000
rect 250866 137944 250871 138000
rect 248860 137942 250871 137944
rect 214097 137939 214163 137942
rect 250805 137939 250871 137942
rect 307569 137866 307635 137869
rect 324313 137866 324379 137869
rect 307569 137864 310132 137866
rect 307569 137808 307574 137864
rect 307630 137808 310132 137864
rect 307569 137806 310132 137808
rect 321908 137864 324379 137866
rect 321908 137808 324318 137864
rect 324374 137808 324379 137864
rect 321908 137806 324379 137808
rect 307569 137803 307635 137806
rect 324313 137803 324379 137806
rect 251265 137594 251331 137597
rect 248860 137592 251331 137594
rect 248860 137536 251270 137592
rect 251326 137536 251331 137592
rect 248860 137534 251331 137536
rect 251265 137531 251331 137534
rect 307477 137458 307543 137461
rect 307477 137456 310132 137458
rect 307477 137400 307482 137456
rect 307538 137400 310132 137456
rect 307477 137398 310132 137400
rect 307477 137395 307543 137398
rect 214649 137322 214715 137325
rect 214649 137320 217212 137322
rect 214649 137264 214654 137320
rect 214710 137264 217212 137320
rect 214649 137262 217212 137264
rect 214649 137259 214715 137262
rect 252461 137050 252527 137053
rect 248860 137048 252527 137050
rect 248860 136992 252466 137048
rect 252522 136992 252527 137048
rect 248860 136990 252527 136992
rect 252461 136987 252527 136990
rect 307661 137050 307727 137053
rect 324497 137050 324563 137053
rect 307661 137048 310132 137050
rect 307661 136992 307666 137048
rect 307722 136992 310132 137048
rect 307661 136990 310132 136992
rect 321908 137048 324563 137050
rect 321908 136992 324502 137048
rect 324558 136992 324563 137048
rect 321908 136990 324563 136992
rect 307661 136987 307727 136990
rect 324497 136987 324563 136990
rect 214005 136642 214071 136645
rect 250529 136642 250595 136645
rect 214005 136640 217212 136642
rect 214005 136584 214010 136640
rect 214066 136584 217212 136640
rect 214005 136582 217212 136584
rect 248860 136640 250595 136642
rect 248860 136584 250534 136640
rect 250590 136584 250595 136640
rect 248860 136582 250595 136584
rect 214005 136579 214071 136582
rect 250529 136579 250595 136582
rect 306925 136642 306991 136645
rect 306925 136640 310132 136642
rect 306925 136584 306930 136640
rect 306986 136584 310132 136640
rect 306925 136582 310132 136584
rect 306925 136579 306991 136582
rect 325877 136370 325943 136373
rect 321908 136368 325943 136370
rect 321908 136312 325882 136368
rect 325938 136312 325943 136368
rect 321908 136310 325943 136312
rect 325877 136307 325943 136310
rect 252461 136234 252527 136237
rect 248860 136232 252527 136234
rect 248860 136176 252466 136232
rect 252522 136176 252527 136232
rect 248860 136174 252527 136176
rect 252461 136171 252527 136174
rect 307477 136234 307543 136237
rect 307477 136232 310132 136234
rect 307477 136176 307482 136232
rect 307538 136176 310132 136232
rect 307477 136174 310132 136176
rect 307477 136171 307543 136174
rect 213913 135962 213979 135965
rect 213913 135960 217212 135962
rect 213913 135904 213918 135960
rect 213974 135904 217212 135960
rect 213913 135902 217212 135904
rect 213913 135899 213979 135902
rect 251725 135690 251791 135693
rect 248860 135688 251791 135690
rect 248860 135632 251730 135688
rect 251786 135632 251791 135688
rect 248860 135630 251791 135632
rect 251725 135627 251791 135630
rect 307661 135690 307727 135693
rect 307661 135688 310132 135690
rect 307661 135632 307666 135688
rect 307722 135632 310132 135688
rect 307661 135630 310132 135632
rect 307661 135627 307727 135630
rect 214557 135282 214623 135285
rect 252093 135282 252159 135285
rect 214557 135280 217212 135282
rect 214557 135224 214562 135280
rect 214618 135224 217212 135280
rect 214557 135222 217212 135224
rect 248860 135280 252159 135282
rect 248860 135224 252098 135280
rect 252154 135224 252159 135280
rect 248860 135222 252159 135224
rect 214557 135219 214623 135222
rect 252093 135219 252159 135222
rect 300158 135220 300164 135284
rect 300228 135282 300234 135284
rect 321878 135282 321938 135524
rect 342294 135282 342300 135284
rect 300228 135222 310132 135282
rect 321878 135222 342300 135282
rect 300228 135220 300234 135222
rect 342294 135220 342300 135222
rect 342364 135220 342370 135284
rect 307477 134874 307543 134877
rect 307477 134872 310132 134874
rect 307477 134816 307482 134872
rect 307538 134816 310132 134872
rect 307477 134814 310132 134816
rect 307477 134811 307543 134814
rect 252461 134738 252527 134741
rect 324313 134738 324379 134741
rect 248860 134736 252527 134738
rect 248860 134680 252466 134736
rect 252522 134680 252527 134736
rect 248860 134678 252527 134680
rect 321908 134736 324379 134738
rect 321908 134680 324318 134736
rect 324374 134680 324379 134736
rect 321908 134678 324379 134680
rect 252461 134675 252527 134678
rect 324313 134675 324379 134678
rect 213913 134602 213979 134605
rect 213913 134600 217212 134602
rect 213913 134544 213918 134600
rect 213974 134544 217212 134600
rect 213913 134542 217212 134544
rect 213913 134539 213979 134542
rect 305729 134466 305795 134469
rect 305729 134464 310132 134466
rect 305729 134408 305734 134464
rect 305790 134408 310132 134464
rect 305729 134406 310132 134408
rect 305729 134403 305795 134406
rect 252277 134330 252343 134333
rect 248860 134328 252343 134330
rect 248860 134272 252282 134328
rect 252338 134272 252343 134328
rect 248860 134270 252343 134272
rect 252277 134267 252343 134270
rect 307661 134058 307727 134061
rect 324497 134058 324563 134061
rect 307661 134056 310132 134058
rect 307661 134000 307666 134056
rect 307722 134000 310132 134056
rect 307661 133998 310132 134000
rect 321908 134056 324563 134058
rect 321908 134000 324502 134056
rect 324558 134000 324563 134056
rect 321908 133998 324563 134000
rect 307661 133995 307727 133998
rect 324497 133995 324563 133998
rect 170254 133860 170260 133924
rect 170324 133922 170330 133924
rect 170324 133862 217212 133922
rect 170324 133860 170330 133862
rect 252461 133786 252527 133789
rect 248860 133784 252527 133786
rect 248860 133728 252466 133784
rect 252522 133728 252527 133784
rect 248860 133726 252527 133728
rect 252461 133723 252527 133726
rect 306925 133650 306991 133653
rect 306925 133648 310132 133650
rect 306925 133592 306930 133648
rect 306986 133592 310132 133648
rect 306925 133590 310132 133592
rect 306925 133587 306991 133590
rect 251265 133378 251331 133381
rect 248860 133376 251331 133378
rect 167678 132772 167684 132836
rect 167748 132834 167754 132836
rect 217182 132834 217242 133348
rect 248860 133320 251270 133376
rect 251326 133320 251331 133376
rect 248860 133318 251331 133320
rect 251265 133315 251331 133318
rect 306557 133242 306623 133245
rect 324313 133242 324379 133245
rect 306557 133240 310132 133242
rect 306557 133184 306562 133240
rect 306618 133184 310132 133240
rect 306557 133182 310132 133184
rect 321908 133240 324379 133242
rect 321908 133184 324318 133240
rect 324374 133184 324379 133240
rect 321908 133182 324379 133184
rect 306557 133179 306623 133182
rect 324313 133179 324379 133182
rect 252369 132834 252435 132837
rect 167748 132774 217242 132834
rect 248860 132832 252435 132834
rect 248860 132776 252374 132832
rect 252430 132776 252435 132832
rect 248860 132774 252435 132776
rect 167748 132772 167754 132774
rect 252369 132771 252435 132774
rect 213913 132698 213979 132701
rect 307661 132698 307727 132701
rect 213913 132696 217212 132698
rect 213913 132640 213918 132696
rect 213974 132640 217212 132696
rect 213913 132638 217212 132640
rect 307661 132696 310132 132698
rect 307661 132640 307666 132696
rect 307722 132640 310132 132696
rect 307661 132638 310132 132640
rect 213913 132635 213979 132638
rect 307661 132635 307727 132638
rect 252185 132426 252251 132429
rect 324313 132426 324379 132429
rect 248860 132424 252251 132426
rect 248860 132368 252190 132424
rect 252246 132368 252251 132424
rect 248860 132366 252251 132368
rect 321908 132424 324379 132426
rect 321908 132368 324318 132424
rect 324374 132368 324379 132424
rect 321908 132366 324379 132368
rect 252185 132363 252251 132366
rect 324313 132363 324379 132366
rect 306925 132290 306991 132293
rect 306925 132288 310132 132290
rect 306925 132232 306930 132288
rect 306986 132232 310132 132288
rect 306925 132230 310132 132232
rect 306925 132227 306991 132230
rect 327574 132154 327580 132156
rect 321878 132094 327580 132154
rect 214833 132018 214899 132021
rect 214833 132016 217212 132018
rect 214833 131960 214838 132016
rect 214894 131960 217212 132016
rect 214833 131958 217212 131960
rect 214833 131955 214899 131958
rect 252277 131882 252343 131885
rect 248860 131880 252343 131882
rect 248860 131824 252282 131880
rect 252338 131824 252343 131880
rect 248860 131822 252343 131824
rect 252277 131819 252343 131822
rect 307661 131882 307727 131885
rect 307661 131880 310132 131882
rect 307661 131824 307666 131880
rect 307722 131824 310132 131880
rect 307661 131822 310132 131824
rect 307661 131819 307727 131822
rect 321878 131716 321938 132094
rect 327574 132092 327580 132094
rect 327644 132092 327650 132156
rect 324405 131746 324471 131749
rect 331254 131746 331260 131748
rect 324405 131744 331260 131746
rect 324405 131688 324410 131744
rect 324466 131688 331260 131744
rect 324405 131686 331260 131688
rect 324405 131683 324471 131686
rect 331254 131684 331260 131686
rect 331324 131684 331330 131748
rect 251725 131474 251791 131477
rect 248860 131472 251791 131474
rect 248860 131416 251730 131472
rect 251786 131416 251791 131472
rect 248860 131414 251791 131416
rect 251725 131411 251791 131414
rect 307385 131474 307451 131477
rect 307385 131472 310132 131474
rect 307385 131416 307390 131472
rect 307446 131416 310132 131472
rect 307385 131414 310132 131416
rect 307385 131411 307451 131414
rect 200070 131278 217212 131338
rect 166206 131140 166212 131204
rect 166276 131202 166282 131204
rect 200070 131202 200130 131278
rect 166276 131142 200130 131202
rect 166276 131140 166282 131142
rect 296670 131006 310132 131066
rect 252461 130930 252527 130933
rect 248860 130928 252527 130930
rect 248860 130872 252466 130928
rect 252522 130872 252527 130928
rect 248860 130870 252527 130872
rect 252461 130867 252527 130870
rect 214005 130658 214071 130661
rect 214005 130656 217212 130658
rect 214005 130600 214010 130656
rect 214066 130600 217212 130656
rect 214005 130598 217212 130600
rect 214005 130595 214071 130598
rect 252369 130522 252435 130525
rect 248860 130520 252435 130522
rect 248860 130464 252374 130520
rect 252430 130464 252435 130520
rect 248860 130462 252435 130464
rect 252369 130459 252435 130462
rect 252277 130114 252343 130117
rect 248860 130112 252343 130114
rect 248860 130056 252282 130112
rect 252338 130056 252343 130112
rect 248860 130054 252343 130056
rect 252277 130051 252343 130054
rect 291694 130052 291700 130116
rect 291764 130114 291770 130116
rect 296670 130114 296730 131006
rect 324405 130930 324471 130933
rect 321908 130928 324471 130930
rect 321908 130872 324410 130928
rect 324466 130872 324471 130928
rect 321908 130870 324471 130872
rect 324405 130867 324471 130870
rect 307109 130658 307175 130661
rect 307109 130656 310132 130658
rect 307109 130600 307114 130656
rect 307170 130600 310132 130656
rect 307109 130598 310132 130600
rect 307109 130595 307175 130598
rect 307661 130250 307727 130253
rect 307661 130248 310132 130250
rect 307661 130192 307666 130248
rect 307722 130192 310132 130248
rect 307661 130190 310132 130192
rect 307661 130187 307727 130190
rect 324313 130114 324379 130117
rect 291764 130054 296730 130114
rect 321908 130112 324379 130114
rect 321908 130056 324318 130112
rect 324374 130056 324379 130112
rect 321908 130054 324379 130056
rect 291764 130052 291770 130054
rect 324313 130051 324379 130054
rect 213913 129978 213979 129981
rect 213913 129976 217212 129978
rect 213913 129920 213918 129976
rect 213974 129920 217212 129976
rect 213913 129918 217212 129920
rect 213913 129915 213979 129918
rect 307293 129842 307359 129845
rect 307293 129840 310132 129842
rect 307293 129784 307298 129840
rect 307354 129784 310132 129840
rect 307293 129782 310132 129784
rect 307293 129779 307359 129782
rect 252461 129570 252527 129573
rect 248860 129568 252527 129570
rect 248860 129512 252466 129568
rect 252522 129512 252527 129568
rect 248860 129510 252527 129512
rect 252461 129507 252527 129510
rect 324313 129434 324379 129437
rect 321908 129432 324379 129434
rect 321908 129376 324318 129432
rect 324374 129376 324379 129432
rect 321908 129374 324379 129376
rect 324313 129371 324379 129374
rect 67541 129298 67607 129301
rect 68142 129298 68816 129304
rect 67541 129296 68816 129298
rect 67541 129240 67546 129296
rect 67602 129244 68816 129296
rect 67602 129240 68202 129244
rect 67541 129238 68202 129240
rect 67541 129235 67607 129238
rect 213913 129298 213979 129301
rect 306741 129298 306807 129301
rect 213913 129296 217212 129298
rect 213913 129240 213918 129296
rect 213974 129240 217212 129296
rect 213913 129238 217212 129240
rect 306741 129296 310132 129298
rect 306741 129240 306746 129296
rect 306802 129240 310132 129296
rect 306741 129238 310132 129240
rect 213913 129235 213979 129238
rect 306741 129235 306807 129238
rect 252369 129162 252435 129165
rect 248860 129160 252435 129162
rect 248860 129104 252374 129160
rect 252430 129104 252435 129160
rect 248860 129102 252435 129104
rect 252369 129099 252435 129102
rect 307661 128890 307727 128893
rect 307661 128888 310132 128890
rect 307661 128832 307666 128888
rect 307722 128832 310132 128888
rect 307661 128830 310132 128832
rect 307661 128827 307727 128830
rect 200070 128694 217212 128754
rect 169150 128556 169156 128620
rect 169220 128618 169226 128620
rect 200070 128618 200130 128694
rect 252277 128618 252343 128621
rect 324405 128618 324471 128621
rect 169220 128558 200130 128618
rect 248860 128616 252343 128618
rect 248860 128560 252282 128616
rect 252338 128560 252343 128616
rect 248860 128558 252343 128560
rect 321908 128616 324471 128618
rect 321908 128560 324410 128616
rect 324466 128560 324471 128616
rect 321908 128558 324471 128560
rect 169220 128556 169226 128558
rect 252277 128555 252343 128558
rect 324405 128555 324471 128558
rect 307293 128482 307359 128485
rect 307293 128480 310132 128482
rect 307293 128424 307298 128480
rect 307354 128424 310132 128480
rect 307293 128422 310132 128424
rect 307293 128419 307359 128422
rect 252461 128210 252527 128213
rect 248860 128208 252527 128210
rect 248860 128152 252466 128208
rect 252522 128152 252527 128208
rect 248860 128150 252527 128152
rect 252461 128147 252527 128150
rect 66161 128074 66227 128077
rect 68142 128074 68816 128080
rect 66161 128072 68816 128074
rect 66161 128016 66166 128072
rect 66222 128020 68816 128072
rect 66222 128016 68202 128020
rect 66161 128014 68202 128016
rect 66161 128011 66227 128014
rect 64781 127122 64847 127125
rect 66161 127122 66227 127125
rect 64781 127120 66227 127122
rect 64781 127064 64786 127120
rect 64842 127064 66166 127120
rect 66222 127064 66227 127120
rect 64781 127062 66227 127064
rect 64781 127059 64847 127062
rect 66161 127059 66227 127062
rect 214005 128074 214071 128077
rect 214005 128072 217212 128074
rect 214005 128016 214010 128072
rect 214066 128016 217212 128072
rect 214005 128014 217212 128016
rect 214005 128011 214071 128014
rect 307150 128012 307156 128076
rect 307220 128074 307226 128076
rect 307220 128014 310132 128074
rect 307220 128012 307226 128014
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 252369 127666 252435 127669
rect 248860 127664 252435 127666
rect 248860 127608 252374 127664
rect 252430 127608 252435 127664
rect 248860 127606 252435 127608
rect 252369 127603 252435 127606
rect 307569 127666 307635 127669
rect 307569 127664 310132 127666
rect 307569 127608 307574 127664
rect 307630 127608 310132 127664
rect 307569 127606 310132 127608
rect 307569 127603 307635 127606
rect 213913 127394 213979 127397
rect 213913 127392 217212 127394
rect 213913 127336 213918 127392
rect 213974 127336 217212 127392
rect 213913 127334 217212 127336
rect 213913 127331 213979 127334
rect 251817 127258 251883 127261
rect 248860 127256 251883 127258
rect 248860 127200 251822 127256
rect 251878 127200 251883 127256
rect 248860 127198 251883 127200
rect 251817 127195 251883 127198
rect 307661 127258 307727 127261
rect 307661 127256 310132 127258
rect 307661 127200 307666 127256
rect 307722 127200 310132 127256
rect 307661 127198 310132 127200
rect 307661 127195 307727 127198
rect 324405 127122 324471 127125
rect 321908 127120 324471 127122
rect 321908 127064 324410 127120
rect 324466 127064 324471 127120
rect 321908 127062 324471 127064
rect 324405 127059 324471 127062
rect 296670 126790 310132 126850
rect 213913 126714 213979 126717
rect 252461 126714 252527 126717
rect 213913 126712 217212 126714
rect 213913 126656 213918 126712
rect 213974 126656 217212 126712
rect 213913 126654 217212 126656
rect 248860 126712 252527 126714
rect 248860 126656 252466 126712
rect 252522 126656 252527 126712
rect 248860 126654 252527 126656
rect 213913 126651 213979 126654
rect 252461 126651 252527 126654
rect 66161 126306 66227 126309
rect 68142 126306 68816 126312
rect 66161 126304 68816 126306
rect 66161 126248 66166 126304
rect 66222 126252 68816 126304
rect 251725 126306 251791 126309
rect 66222 126248 68202 126252
rect 66161 126246 68202 126248
rect 66161 126243 66227 126246
rect 248860 126304 251791 126306
rect 248860 126248 251730 126304
rect 251786 126248 251791 126304
rect 248860 126246 251791 126248
rect 251725 126243 251791 126246
rect 214741 126034 214807 126037
rect 214741 126032 217212 126034
rect 214741 125976 214746 126032
rect 214802 125976 217212 126032
rect 214741 125974 217212 125976
rect 214741 125971 214807 125974
rect 293166 125836 293172 125900
rect 293236 125898 293242 125900
rect 296670 125898 296730 126790
rect 306557 126442 306623 126445
rect 306557 126440 310132 126442
rect 306557 126384 306562 126440
rect 306618 126384 310132 126440
rect 306557 126382 310132 126384
rect 306557 126379 306623 126382
rect 324313 126306 324379 126309
rect 321908 126304 324379 126306
rect 321908 126248 324318 126304
rect 324374 126248 324379 126304
rect 321908 126246 324379 126248
rect 324313 126243 324379 126246
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 293236 125838 296730 125898
rect 306925 125898 306991 125901
rect 306925 125896 310132 125898
rect 306925 125840 306930 125896
rect 306986 125840 310132 125896
rect 583520 125884 584960 125974
rect 306925 125838 310132 125840
rect 293236 125836 293242 125838
rect 306925 125835 306991 125838
rect 252185 125762 252251 125765
rect 248860 125760 252251 125762
rect 248860 125704 252190 125760
rect 252246 125704 252251 125760
rect 248860 125702 252251 125704
rect 252185 125699 252251 125702
rect 306925 125490 306991 125493
rect 324497 125490 324563 125493
rect 306925 125488 310132 125490
rect 306925 125432 306930 125488
rect 306986 125432 310132 125488
rect 306925 125430 310132 125432
rect 321908 125488 324563 125490
rect 321908 125432 324502 125488
rect 324558 125432 324563 125488
rect 321908 125430 324563 125432
rect 306925 125427 306991 125430
rect 324497 125427 324563 125430
rect 214005 125354 214071 125357
rect 252461 125354 252527 125357
rect 214005 125352 217212 125354
rect 214005 125296 214010 125352
rect 214066 125296 217212 125352
rect 214005 125294 217212 125296
rect 248860 125352 252527 125354
rect 248860 125296 252466 125352
rect 252522 125296 252527 125352
rect 248860 125294 252527 125296
rect 214005 125291 214071 125294
rect 252461 125291 252527 125294
rect 66161 125218 66227 125221
rect 68142 125218 68816 125224
rect 66161 125216 68816 125218
rect 66161 125160 66166 125216
rect 66222 125164 68816 125216
rect 66222 125160 68202 125164
rect 66161 125158 68202 125160
rect 66161 125155 66227 125158
rect -960 123572 480 123812
rect 307477 125082 307543 125085
rect 307477 125080 310132 125082
rect 307477 125024 307482 125080
rect 307538 125024 310132 125080
rect 307477 125022 310132 125024
rect 307477 125019 307543 125022
rect 252093 124810 252159 124813
rect 325601 124810 325667 124813
rect 248860 124808 252159 124810
rect 248860 124752 252098 124808
rect 252154 124752 252159 124808
rect 248860 124750 252159 124752
rect 321908 124808 325667 124810
rect 321908 124752 325606 124808
rect 325662 124752 325667 124808
rect 321908 124750 325667 124752
rect 252093 124747 252159 124750
rect 325601 124747 325667 124750
rect 213913 124674 213979 124677
rect 305637 124674 305703 124677
rect 213913 124672 217212 124674
rect 213913 124616 213918 124672
rect 213974 124616 217212 124672
rect 213913 124614 217212 124616
rect 305637 124672 310132 124674
rect 305637 124616 305642 124672
rect 305698 124616 310132 124672
rect 305637 124614 310132 124616
rect 213913 124611 213979 124614
rect 305637 124611 305703 124614
rect 252461 124402 252527 124405
rect 248860 124400 252527 124402
rect 248860 124344 252466 124400
rect 252522 124344 252527 124400
rect 248860 124342 252527 124344
rect 252461 124339 252527 124342
rect 307661 124266 307727 124269
rect 307661 124264 310132 124266
rect 307661 124208 307666 124264
rect 307722 124208 310132 124264
rect 307661 124206 310132 124208
rect 307661 124203 307727 124206
rect 214005 124130 214071 124133
rect 214005 124128 217212 124130
rect 214005 124072 214010 124128
rect 214066 124072 217212 124128
rect 214005 124070 217212 124072
rect 214005 124067 214071 124070
rect 251541 123994 251607 123997
rect 248860 123992 251607 123994
rect 248860 123936 251546 123992
rect 251602 123936 251607 123992
rect 248860 123934 251607 123936
rect 251541 123931 251607 123934
rect 307569 123858 307635 123861
rect 307569 123856 310132 123858
rect 307569 123800 307574 123856
rect 307630 123800 310132 123856
rect 307569 123798 310132 123800
rect 307569 123795 307635 123798
rect 67449 123586 67515 123589
rect 68142 123586 68816 123592
rect 67449 123584 68816 123586
rect 67449 123528 67454 123584
rect 67510 123532 68816 123584
rect 67510 123528 68202 123532
rect 67449 123526 68202 123528
rect 67449 123523 67515 123526
rect 213913 123450 213979 123453
rect 252461 123450 252527 123453
rect 213913 123448 217212 123450
rect 213913 123392 213918 123448
rect 213974 123392 217212 123448
rect 213913 123390 217212 123392
rect 248860 123448 252527 123450
rect 248860 123392 252466 123448
rect 252522 123392 252527 123448
rect 248860 123390 252527 123392
rect 213913 123387 213979 123390
rect 252461 123387 252527 123390
rect 307661 123450 307727 123453
rect 307661 123448 310132 123450
rect 307661 123392 307666 123448
rect 307722 123392 310132 123448
rect 307661 123390 310132 123392
rect 307661 123387 307727 123390
rect 321878 123314 321938 123964
rect 332726 123314 332732 123316
rect 321878 123254 332732 123314
rect 332726 123252 332732 123254
rect 332796 123252 332802 123316
rect 324313 123178 324379 123181
rect 321908 123176 324379 123178
rect 321908 123120 324318 123176
rect 324374 123120 324379 123176
rect 321908 123118 324379 123120
rect 324313 123115 324379 123118
rect 251265 123042 251331 123045
rect 248860 123040 251331 123042
rect 248860 122984 251270 123040
rect 251326 122984 251331 123040
rect 248860 122982 251331 122984
rect 251265 122979 251331 122982
rect 307477 123042 307543 123045
rect 307477 123040 310132 123042
rect 307477 122984 307482 123040
rect 307538 122984 310132 123040
rect 307477 122982 310132 122984
rect 307477 122979 307543 122982
rect 214005 122770 214071 122773
rect 214005 122768 217212 122770
rect 214005 122712 214010 122768
rect 214066 122712 217212 122768
rect 214005 122710 217212 122712
rect 214005 122707 214071 122710
rect 66069 122634 66135 122637
rect 68142 122634 68816 122640
rect 66069 122632 68816 122634
rect 66069 122576 66074 122632
rect 66130 122580 68816 122632
rect 66130 122576 68202 122580
rect 66069 122574 68202 122576
rect 66069 122571 66135 122574
rect 252461 122498 252527 122501
rect 248860 122496 252527 122498
rect 248860 122440 252466 122496
rect 252522 122440 252527 122496
rect 248860 122438 252527 122440
rect 252461 122435 252527 122438
rect 307477 122498 307543 122501
rect 324313 122498 324379 122501
rect 307477 122496 310132 122498
rect 307477 122440 307482 122496
rect 307538 122440 310132 122496
rect 307477 122438 310132 122440
rect 321908 122496 324379 122498
rect 321908 122440 324318 122496
rect 324374 122440 324379 122496
rect 321908 122438 324379 122440
rect 307477 122435 307543 122438
rect 324313 122435 324379 122438
rect 213913 122090 213979 122093
rect 251725 122090 251791 122093
rect 213913 122088 217212 122090
rect 213913 122032 213918 122088
rect 213974 122032 217212 122088
rect 213913 122030 217212 122032
rect 248860 122088 251791 122090
rect 248860 122032 251730 122088
rect 251786 122032 251791 122088
rect 248860 122030 251791 122032
rect 213913 122027 213979 122030
rect 251725 122027 251791 122030
rect 307661 122090 307727 122093
rect 307661 122088 310132 122090
rect 307661 122032 307666 122088
rect 307722 122032 310132 122088
rect 307661 122030 310132 122032
rect 307661 122027 307727 122030
rect 306925 121682 306991 121685
rect 324405 121682 324471 121685
rect 306925 121680 310132 121682
rect 306925 121624 306930 121680
rect 306986 121624 310132 121680
rect 306925 121622 310132 121624
rect 321908 121680 324471 121682
rect 321908 121624 324410 121680
rect 324466 121624 324471 121680
rect 321908 121622 324471 121624
rect 306925 121619 306991 121622
rect 324405 121619 324471 121622
rect 252369 121546 252435 121549
rect 248860 121544 252435 121546
rect 248860 121488 252374 121544
rect 252430 121488 252435 121544
rect 248860 121486 252435 121488
rect 252369 121483 252435 121486
rect 213269 121410 213335 121413
rect 213269 121408 217212 121410
rect 213269 121352 213274 121408
rect 213330 121352 217212 121408
rect 213269 121350 217212 121352
rect 213269 121347 213335 121350
rect 306741 121274 306807 121277
rect 306741 121272 310132 121274
rect 306741 121216 306746 121272
rect 306802 121216 310132 121272
rect 306741 121214 310132 121216
rect 306741 121211 306807 121214
rect 252461 121138 252527 121141
rect 248860 121136 252527 121138
rect 248860 121080 252466 121136
rect 252522 121080 252527 121136
rect 248860 121078 252527 121080
rect 252461 121075 252527 121078
rect 67357 120866 67423 120869
rect 68142 120866 68816 120872
rect 67357 120864 68816 120866
rect 67357 120808 67362 120864
rect 67418 120812 68816 120864
rect 67418 120808 68202 120812
rect 67357 120806 68202 120808
rect 67357 120803 67423 120806
rect 307477 120866 307543 120869
rect 324313 120866 324379 120869
rect 307477 120864 310132 120866
rect 307477 120808 307482 120864
rect 307538 120808 310132 120864
rect 307477 120806 310132 120808
rect 321908 120864 324379 120866
rect 321908 120808 324318 120864
rect 324374 120808 324379 120864
rect 321908 120806 324379 120808
rect 307477 120803 307543 120806
rect 324313 120803 324379 120806
rect 213913 120730 213979 120733
rect 213913 120728 217212 120730
rect 213913 120672 213918 120728
rect 213974 120672 217212 120728
rect 213913 120670 217212 120672
rect 213913 120667 213979 120670
rect 251725 120594 251791 120597
rect 248860 120592 251791 120594
rect 248860 120536 251730 120592
rect 251786 120536 251791 120592
rect 248860 120534 251791 120536
rect 251725 120531 251791 120534
rect 307661 120458 307727 120461
rect 307661 120456 310132 120458
rect 307661 120400 307666 120456
rect 307722 120400 310132 120456
rect 307661 120398 310132 120400
rect 307661 120395 307727 120398
rect 252369 120186 252435 120189
rect 324405 120186 324471 120189
rect 248860 120184 252435 120186
rect 248860 120128 252374 120184
rect 252430 120128 252435 120184
rect 248860 120126 252435 120128
rect 321908 120184 324471 120186
rect 321908 120128 324410 120184
rect 324466 120128 324471 120184
rect 321908 120126 324471 120128
rect 252369 120123 252435 120126
rect 324405 120123 324471 120126
rect 214097 120050 214163 120053
rect 306925 120050 306991 120053
rect 214097 120048 217212 120050
rect 214097 119992 214102 120048
rect 214158 119992 217212 120048
rect 214097 119990 217212 119992
rect 306925 120048 310132 120050
rect 306925 119992 306930 120048
rect 306986 119992 310132 120048
rect 306925 119990 310132 119992
rect 214097 119987 214163 119990
rect 306925 119987 306991 119990
rect 252277 119642 252343 119645
rect 248860 119640 252343 119642
rect 248860 119584 252282 119640
rect 252338 119584 252343 119640
rect 248860 119582 252343 119584
rect 252277 119579 252343 119582
rect 306557 119642 306623 119645
rect 306557 119640 310132 119642
rect 306557 119584 306562 119640
rect 306618 119584 310132 119640
rect 306557 119582 310132 119584
rect 306557 119579 306623 119582
rect 214005 119506 214071 119509
rect 214005 119504 217212 119506
rect 214005 119448 214010 119504
rect 214066 119448 217212 119504
rect 214005 119446 217212 119448
rect 214005 119443 214071 119446
rect 324313 119370 324379 119373
rect 321908 119368 324379 119370
rect 321908 119312 324318 119368
rect 324374 119312 324379 119368
rect 321908 119310 324379 119312
rect 324313 119307 324379 119310
rect 252185 119234 252251 119237
rect 248860 119232 252251 119234
rect 248860 119176 252190 119232
rect 252246 119176 252251 119232
rect 248860 119174 252251 119176
rect 252185 119171 252251 119174
rect 307661 119098 307727 119101
rect 307661 119096 310132 119098
rect 307661 119040 307666 119096
rect 307722 119040 310132 119096
rect 307661 119038 310132 119040
rect 307661 119035 307727 119038
rect 213913 118826 213979 118829
rect 251449 118826 251515 118829
rect 213913 118824 217212 118826
rect 213913 118768 213918 118824
rect 213974 118768 217212 118824
rect 213913 118766 217212 118768
rect 248860 118824 251515 118826
rect 248860 118768 251454 118824
rect 251510 118768 251515 118824
rect 248860 118766 251515 118768
rect 213913 118763 213979 118766
rect 251449 118763 251515 118766
rect 307569 118690 307635 118693
rect 307569 118688 310132 118690
rect 307569 118632 307574 118688
rect 307630 118632 310132 118688
rect 307569 118630 310132 118632
rect 307569 118627 307635 118630
rect 324313 118554 324379 118557
rect 321908 118552 324379 118554
rect 321908 118496 324318 118552
rect 324374 118496 324379 118552
rect 321908 118494 324379 118496
rect 324313 118491 324379 118494
rect 252461 118282 252527 118285
rect 248860 118280 252527 118282
rect 248860 118224 252466 118280
rect 252522 118224 252527 118280
rect 248860 118222 252527 118224
rect 252461 118219 252527 118222
rect 306557 118282 306623 118285
rect 306557 118280 310132 118282
rect 306557 118224 306562 118280
rect 306618 118224 310132 118280
rect 306557 118222 310132 118224
rect 306557 118219 306623 118222
rect 214005 118146 214071 118149
rect 214005 118144 217212 118146
rect 214005 118088 214010 118144
rect 214066 118088 217212 118144
rect 214005 118086 217212 118088
rect 214005 118083 214071 118086
rect 251725 117874 251791 117877
rect 248860 117872 251791 117874
rect 248860 117816 251730 117872
rect 251786 117816 251791 117872
rect 248860 117814 251791 117816
rect 251725 117811 251791 117814
rect 307661 117874 307727 117877
rect 324405 117874 324471 117877
rect 307661 117872 310132 117874
rect 307661 117816 307666 117872
rect 307722 117816 310132 117872
rect 307661 117814 310132 117816
rect 321908 117872 324471 117874
rect 321908 117816 324410 117872
rect 324466 117816 324471 117872
rect 321908 117814 324471 117816
rect 307661 117811 307727 117814
rect 324405 117811 324471 117814
rect 295926 117540 295932 117604
rect 295996 117602 296002 117604
rect 295996 117542 296730 117602
rect 295996 117540 296002 117542
rect 213913 117466 213979 117469
rect 296670 117466 296730 117542
rect 213913 117464 217212 117466
rect 213913 117408 213918 117464
rect 213974 117408 217212 117464
rect 213913 117406 217212 117408
rect 296670 117406 310132 117466
rect 213913 117403 213979 117406
rect 252277 117330 252343 117333
rect 248860 117328 252343 117330
rect 248860 117272 252282 117328
rect 252338 117272 252343 117328
rect 248860 117270 252343 117272
rect 252277 117267 252343 117270
rect 306741 117058 306807 117061
rect 306741 117056 310132 117058
rect 306741 117000 306746 117056
rect 306802 117000 310132 117056
rect 306741 116998 310132 117000
rect 306741 116995 306807 116998
rect 251265 116922 251331 116925
rect 248860 116920 251331 116922
rect 248860 116864 251270 116920
rect 251326 116864 251331 116920
rect 248860 116862 251331 116864
rect 251265 116859 251331 116862
rect 214005 116786 214071 116789
rect 214005 116784 217212 116786
rect 214005 116728 214010 116784
rect 214066 116728 217212 116784
rect 214005 116726 217212 116728
rect 214005 116723 214071 116726
rect 307569 116650 307635 116653
rect 307569 116648 310132 116650
rect 307569 116592 307574 116648
rect 307630 116592 310132 116648
rect 307569 116590 310132 116592
rect 307569 116587 307635 116590
rect 321878 116514 321938 117028
rect 323485 116514 323551 116517
rect 321878 116512 323551 116514
rect 321878 116456 323490 116512
rect 323546 116456 323551 116512
rect 321878 116454 323551 116456
rect 323485 116451 323551 116454
rect 252461 116378 252527 116381
rect 248860 116376 252527 116378
rect 248860 116320 252466 116376
rect 252522 116320 252527 116376
rect 248860 116318 252527 116320
rect 252461 116315 252527 116318
rect 307661 116242 307727 116245
rect 307661 116240 310132 116242
rect 307661 116184 307666 116240
rect 307722 116184 310132 116240
rect 307661 116182 310132 116184
rect 307661 116179 307727 116182
rect 213913 116106 213979 116109
rect 321878 116106 321938 116348
rect 335670 116106 335676 116108
rect 213913 116104 217212 116106
rect 213913 116048 213918 116104
rect 213974 116048 217212 116104
rect 213913 116046 217212 116048
rect 321878 116046 335676 116106
rect 213913 116043 213979 116046
rect 335670 116044 335676 116046
rect 335740 116044 335746 116108
rect 251909 115970 251975 115973
rect 248860 115968 251975 115970
rect 248860 115912 251914 115968
rect 251970 115912 251975 115968
rect 248860 115910 251975 115912
rect 251909 115907 251975 115910
rect 323485 115970 323551 115973
rect 338246 115970 338252 115972
rect 323485 115968 338252 115970
rect 323485 115912 323490 115968
rect 323546 115912 338252 115968
rect 323485 115910 338252 115912
rect 323485 115907 323551 115910
rect 338246 115908 338252 115910
rect 338316 115908 338322 115972
rect 306741 115698 306807 115701
rect 306741 115696 310132 115698
rect 306741 115640 306746 115696
rect 306802 115640 310132 115696
rect 306741 115638 310132 115640
rect 306741 115635 306807 115638
rect 324313 115562 324379 115565
rect 321908 115560 324379 115562
rect 321908 115504 324318 115560
rect 324374 115504 324379 115560
rect 321908 115502 324379 115504
rect 324313 115499 324379 115502
rect 214005 115426 214071 115429
rect 251541 115426 251607 115429
rect 214005 115424 217212 115426
rect 214005 115368 214010 115424
rect 214066 115368 217212 115424
rect 214005 115366 217212 115368
rect 248860 115424 251607 115426
rect 248860 115368 251546 115424
rect 251602 115368 251607 115424
rect 248860 115366 251607 115368
rect 214005 115363 214071 115366
rect 251541 115363 251607 115366
rect 307569 115290 307635 115293
rect 307569 115288 310132 115290
rect 307569 115232 307574 115288
rect 307630 115232 310132 115288
rect 307569 115230 310132 115232
rect 307569 115227 307635 115230
rect 251950 115092 251956 115156
rect 252020 115154 252026 115156
rect 304349 115154 304415 115157
rect 252020 115152 304415 115154
rect 252020 115096 304354 115152
rect 304410 115096 304415 115152
rect 252020 115094 304415 115096
rect 252020 115092 252026 115094
rect 304349 115091 304415 115094
rect 251173 115018 251239 115021
rect 248860 115016 251239 115018
rect 248860 114960 251178 115016
rect 251234 114960 251239 115016
rect 248860 114958 251239 114960
rect 251173 114955 251239 114958
rect 213913 114882 213979 114885
rect 307661 114882 307727 114885
rect 213913 114880 217212 114882
rect 213913 114824 213918 114880
rect 213974 114824 217212 114880
rect 213913 114822 217212 114824
rect 307661 114880 310132 114882
rect 307661 114824 307666 114880
rect 307722 114824 310132 114880
rect 307661 114822 310132 114824
rect 213913 114819 213979 114822
rect 307661 114819 307727 114822
rect 324405 114746 324471 114749
rect 321908 114744 324471 114746
rect 321908 114688 324410 114744
rect 324466 114688 324471 114744
rect 321908 114686 324471 114688
rect 324405 114683 324471 114686
rect 252461 114474 252527 114477
rect 248860 114472 252527 114474
rect 248860 114416 252466 114472
rect 252522 114416 252527 114472
rect 248860 114414 252527 114416
rect 252461 114411 252527 114414
rect 296670 114414 310132 114474
rect 214005 114202 214071 114205
rect 214005 114200 217212 114202
rect 214005 114144 214010 114200
rect 214066 114144 217212 114200
rect 214005 114142 217212 114144
rect 214005 114139 214071 114142
rect 252369 114066 252435 114069
rect 248860 114064 252435 114066
rect 248860 114008 252374 114064
rect 252430 114008 252435 114064
rect 248860 114006 252435 114008
rect 252369 114003 252435 114006
rect 213913 113522 213979 113525
rect 252461 113522 252527 113525
rect 213913 113520 217212 113522
rect 213913 113464 213918 113520
rect 213974 113464 217212 113520
rect 213913 113462 217212 113464
rect 248860 113520 252527 113522
rect 248860 113464 252466 113520
rect 252522 113464 252527 113520
rect 248860 113462 252527 113464
rect 213913 113459 213979 113462
rect 252461 113459 252527 113462
rect 275134 113460 275140 113524
rect 275204 113522 275210 113524
rect 296670 113522 296730 114414
rect 307017 114066 307083 114069
rect 324313 114066 324379 114069
rect 307017 114064 310132 114066
rect 307017 114008 307022 114064
rect 307078 114008 310132 114064
rect 307017 114006 310132 114008
rect 321908 114064 324379 114066
rect 321908 114008 324318 114064
rect 324374 114008 324379 114064
rect 321908 114006 324379 114008
rect 307017 114003 307083 114006
rect 324313 114003 324379 114006
rect 307569 113658 307635 113661
rect 307569 113656 310132 113658
rect 307569 113600 307574 113656
rect 307630 113600 310132 113656
rect 307569 113598 310132 113600
rect 307569 113595 307635 113598
rect 275204 113462 296730 113522
rect 275204 113460 275210 113462
rect 307661 113250 307727 113253
rect 324405 113250 324471 113253
rect 307661 113248 310132 113250
rect 307661 113192 307666 113248
rect 307722 113192 310132 113248
rect 307661 113190 310132 113192
rect 321908 113248 324471 113250
rect 321908 113192 324410 113248
rect 324466 113192 324471 113248
rect 321908 113190 324471 113192
rect 307661 113187 307727 113190
rect 324405 113187 324471 113190
rect 251766 113114 251772 113116
rect 248860 113054 251772 113114
rect 251766 113052 251772 113054
rect 251836 113052 251842 113116
rect 214005 112842 214071 112845
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 214005 112840 217212 112842
rect 214005 112784 214010 112840
rect 214066 112784 217212 112840
rect 214005 112782 217212 112784
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 214005 112779 214071 112782
rect 579797 112779 579863 112782
rect 251725 112706 251791 112709
rect 248860 112704 251791 112706
rect 248860 112648 251730 112704
rect 251786 112648 251791 112704
rect 248860 112646 251791 112648
rect 251725 112643 251791 112646
rect 307477 112706 307543 112709
rect 307477 112704 310132 112706
rect 307477 112648 307482 112704
rect 307538 112648 310132 112704
rect 583520 112692 584960 112782
rect 307477 112646 310132 112648
rect 307477 112643 307543 112646
rect 324313 112434 324379 112437
rect 321908 112432 324379 112434
rect 321908 112376 324318 112432
rect 324374 112376 324379 112432
rect 321908 112374 324379 112376
rect 324313 112371 324379 112374
rect 307569 112298 307635 112301
rect 307569 112296 310132 112298
rect 307569 112240 307574 112296
rect 307630 112240 310132 112296
rect 307569 112238 310132 112240
rect 307569 112235 307635 112238
rect 213913 112162 213979 112165
rect 252093 112162 252159 112165
rect 213913 112160 217212 112162
rect 213913 112104 213918 112160
rect 213974 112104 217212 112160
rect 213913 112102 217212 112104
rect 248860 112160 252159 112162
rect 248860 112104 252098 112160
rect 252154 112104 252159 112160
rect 248860 112102 252159 112104
rect 213913 112099 213979 112102
rect 252093 112099 252159 112102
rect 307661 111890 307727 111893
rect 307661 111888 310132 111890
rect 307661 111832 307666 111888
rect 307722 111832 310132 111888
rect 307661 111830 310132 111832
rect 307661 111827 307727 111830
rect 167913 111754 167979 111757
rect 252001 111754 252067 111757
rect 324313 111754 324379 111757
rect 164694 111752 167979 111754
rect 164694 111696 167918 111752
rect 167974 111696 167979 111752
rect 164694 111694 167979 111696
rect 248860 111752 252067 111754
rect 248860 111696 252006 111752
rect 252062 111696 252067 111752
rect 248860 111694 252067 111696
rect 321908 111752 324379 111754
rect 321908 111696 324318 111752
rect 324374 111696 324379 111752
rect 321908 111694 324379 111696
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 167913 111691 167979 111694
rect 252001 111691 252067 111694
rect 324313 111691 324379 111694
rect 214005 111482 214071 111485
rect 307477 111482 307543 111485
rect 214005 111480 217212 111482
rect 214005 111424 214010 111480
rect 214066 111424 217212 111480
rect 214005 111422 217212 111424
rect 307477 111480 310132 111482
rect 307477 111424 307482 111480
rect 307538 111424 310132 111480
rect 307477 111422 310132 111424
rect 214005 111419 214071 111422
rect 307477 111419 307543 111422
rect 251633 111210 251699 111213
rect 248860 111208 251699 111210
rect 248860 111152 251638 111208
rect 251694 111152 251699 111208
rect 248860 111150 251699 111152
rect 251633 111147 251699 111150
rect 307661 111074 307727 111077
rect 307661 111072 310132 111074
rect 307661 111016 307666 111072
rect 307722 111016 310132 111072
rect 307661 111014 310132 111016
rect 307661 111011 307727 111014
rect 324405 110938 324471 110941
rect 321908 110936 324471 110938
rect 321908 110880 324410 110936
rect 324466 110880 324471 110936
rect 321908 110878 324471 110880
rect 324405 110875 324471 110878
rect 213913 110802 213979 110805
rect 252093 110802 252159 110805
rect 213913 110800 217212 110802
rect 213913 110744 213918 110800
rect 213974 110744 217212 110800
rect 213913 110742 217212 110744
rect 248860 110800 252159 110802
rect 248860 110744 252098 110800
rect 252154 110744 252159 110800
rect 248860 110742 252159 110744
rect 213913 110739 213979 110742
rect 252093 110739 252159 110742
rect 307569 110666 307635 110669
rect 307569 110664 310132 110666
rect 307569 110608 307574 110664
rect 307630 110608 310132 110664
rect 307569 110606 310132 110608
rect 307569 110603 307635 110606
rect 214005 110258 214071 110261
rect 251541 110258 251607 110261
rect 214005 110256 217212 110258
rect 214005 110200 214010 110256
rect 214066 110200 217212 110256
rect 214005 110198 217212 110200
rect 248860 110256 251607 110258
rect 248860 110200 251546 110256
rect 251602 110200 251607 110256
rect 248860 110198 251607 110200
rect 214005 110195 214071 110198
rect 251541 110195 251607 110198
rect 307477 110258 307543 110261
rect 307477 110256 310132 110258
rect 307477 110200 307482 110256
rect 307538 110200 310132 110256
rect 307477 110198 310132 110200
rect 307477 110195 307543 110198
rect 168097 110122 168163 110125
rect 324313 110122 324379 110125
rect 164694 110120 168163 110122
rect 164694 110064 168102 110120
rect 168158 110064 168163 110120
rect 164694 110062 168163 110064
rect 321908 110120 324379 110122
rect 321908 110064 324318 110120
rect 324374 110064 324379 110120
rect 321908 110062 324379 110064
rect 168097 110059 168163 110062
rect 324313 110059 324379 110062
rect 252461 109850 252527 109853
rect 248860 109848 252527 109850
rect 248860 109792 252466 109848
rect 252522 109792 252527 109848
rect 248860 109790 252527 109792
rect 252461 109787 252527 109790
rect 307569 109850 307635 109853
rect 307569 109848 310132 109850
rect 307569 109792 307574 109848
rect 307630 109792 310132 109848
rect 307569 109790 310132 109792
rect 307569 109787 307635 109790
rect 213913 109578 213979 109581
rect 213913 109576 217212 109578
rect 213913 109520 213918 109576
rect 213974 109520 217212 109576
rect 213913 109518 217212 109520
rect 213913 109515 213979 109518
rect 252093 109306 252159 109309
rect 248860 109304 252159 109306
rect 248860 109248 252098 109304
rect 252154 109248 252159 109304
rect 248860 109246 252159 109248
rect 252093 109243 252159 109246
rect 307661 109306 307727 109309
rect 307661 109304 310132 109306
rect 307661 109248 307666 109304
rect 307722 109248 310132 109304
rect 307661 109246 310132 109248
rect 307661 109243 307727 109246
rect 321878 109170 321938 109412
rect 336774 109170 336780 109172
rect 321878 109110 336780 109170
rect 336774 109108 336780 109110
rect 336844 109108 336850 109172
rect 214005 108898 214071 108901
rect 252461 108898 252527 108901
rect 214005 108896 217212 108898
rect 214005 108840 214010 108896
rect 214066 108840 217212 108896
rect 214005 108838 217212 108840
rect 248860 108896 252527 108898
rect 248860 108840 252466 108896
rect 252522 108840 252527 108896
rect 248860 108838 252527 108840
rect 214005 108835 214071 108838
rect 252461 108835 252527 108838
rect 307477 108898 307543 108901
rect 307477 108896 310132 108898
rect 307477 108840 307482 108896
rect 307538 108840 310132 108896
rect 307477 108838 310132 108840
rect 307477 108835 307543 108838
rect 167913 108762 167979 108765
rect 164694 108760 167979 108762
rect 164694 108704 167918 108760
rect 167974 108704 167979 108760
rect 164694 108702 167979 108704
rect 167913 108699 167979 108702
rect 323117 108626 323183 108629
rect 321908 108624 323183 108626
rect 321908 108568 323122 108624
rect 323178 108568 323183 108624
rect 321908 108566 323183 108568
rect 323117 108563 323183 108566
rect 307569 108490 307635 108493
rect 307569 108488 310132 108490
rect 307569 108432 307574 108488
rect 307630 108432 310132 108488
rect 307569 108430 310132 108432
rect 307569 108427 307635 108430
rect 252185 108354 252251 108357
rect 248860 108352 252251 108354
rect 248860 108296 252190 108352
rect 252246 108296 252251 108352
rect 248860 108294 252251 108296
rect 252185 108291 252251 108294
rect 213913 108218 213979 108221
rect 213913 108216 217212 108218
rect 213913 108160 213918 108216
rect 213974 108160 217212 108216
rect 213913 108158 217212 108160
rect 213913 108155 213979 108158
rect 306925 108082 306991 108085
rect 306925 108080 310132 108082
rect 306925 108024 306930 108080
rect 306986 108024 310132 108080
rect 306925 108022 310132 108024
rect 306925 108019 306991 108022
rect 252001 107946 252067 107949
rect 248860 107944 252067 107946
rect 248860 107888 252006 107944
rect 252062 107888 252067 107944
rect 248860 107886 252067 107888
rect 252001 107883 252067 107886
rect 305821 107810 305887 107813
rect 307477 107810 307543 107813
rect 305821 107808 307543 107810
rect 305821 107752 305826 107808
rect 305882 107752 307482 107808
rect 307538 107752 307543 107808
rect 305821 107750 307543 107752
rect 305821 107747 305887 107750
rect 307477 107747 307543 107750
rect 307661 107674 307727 107677
rect 307661 107672 310132 107674
rect 307661 107616 307666 107672
rect 307722 107616 310132 107672
rect 307661 107614 310132 107616
rect 307661 107611 307727 107614
rect 321694 107541 321754 107780
rect 214005 107538 214071 107541
rect 252461 107538 252527 107541
rect 214005 107536 217212 107538
rect 214005 107480 214010 107536
rect 214066 107480 217212 107536
rect 214005 107478 217212 107480
rect 248860 107536 252527 107538
rect 248860 107480 252466 107536
rect 252522 107480 252527 107536
rect 248860 107478 252527 107480
rect 214005 107475 214071 107478
rect 252461 107475 252527 107478
rect 321645 107536 321754 107541
rect 321645 107480 321650 107536
rect 321706 107480 321754 107536
rect 321645 107478 321754 107480
rect 321645 107475 321711 107478
rect 307477 107266 307543 107269
rect 307477 107264 310132 107266
rect 307477 107208 307482 107264
rect 307538 107208 310132 107264
rect 307477 107206 310132 107208
rect 307477 107203 307543 107206
rect 323025 107130 323091 107133
rect 321908 107128 323091 107130
rect 321908 107072 323030 107128
rect 323086 107072 323091 107128
rect 321908 107070 323091 107072
rect 323025 107067 323091 107070
rect 251817 106994 251883 106997
rect 248860 106992 251883 106994
rect 248860 106936 251822 106992
rect 251878 106936 251883 106992
rect 248860 106934 251883 106936
rect 251817 106931 251883 106934
rect 213913 106858 213979 106861
rect 307569 106858 307635 106861
rect 213913 106856 217212 106858
rect 213913 106800 213918 106856
rect 213974 106800 217212 106856
rect 213913 106798 217212 106800
rect 307569 106856 310132 106858
rect 307569 106800 307574 106856
rect 307630 106800 310132 106856
rect 307569 106798 310132 106800
rect 213913 106795 213979 106798
rect 307569 106795 307635 106798
rect 252093 106586 252159 106589
rect 248860 106584 252159 106586
rect 248860 106528 252098 106584
rect 252154 106528 252159 106584
rect 248860 106526 252159 106528
rect 252093 106523 252159 106526
rect 307661 106450 307727 106453
rect 307661 106448 310132 106450
rect 307661 106392 307666 106448
rect 307722 106392 310132 106448
rect 307661 106390 310132 106392
rect 307661 106387 307727 106390
rect 322933 106314 322999 106317
rect 321908 106312 322999 106314
rect 321908 106256 322938 106312
rect 322994 106256 322999 106312
rect 321908 106254 322999 106256
rect 322933 106251 322999 106254
rect 214097 106178 214163 106181
rect 214097 106176 217212 106178
rect 214097 106120 214102 106176
rect 214158 106120 217212 106176
rect 214097 106118 217212 106120
rect 214097 106115 214163 106118
rect 252001 106042 252067 106045
rect 321553 106042 321619 106045
rect 248860 106040 252067 106042
rect 248860 105984 252006 106040
rect 252062 105984 252067 106040
rect 248860 105982 252067 105984
rect 252001 105979 252067 105982
rect 321510 106040 321619 106042
rect 321510 105984 321558 106040
rect 321614 105984 321619 106040
rect 321510 105979 321619 105984
rect 307661 105906 307727 105909
rect 307661 105904 310132 105906
rect 307661 105848 307666 105904
rect 307722 105848 310132 105904
rect 307661 105846 310132 105848
rect 307661 105843 307727 105846
rect 214005 105634 214071 105637
rect 252461 105634 252527 105637
rect 214005 105632 217212 105634
rect 214005 105576 214010 105632
rect 214066 105576 217212 105632
rect 214005 105574 217212 105576
rect 248860 105632 252527 105634
rect 248860 105576 252466 105632
rect 252522 105576 252527 105632
rect 248860 105574 252527 105576
rect 214005 105571 214071 105574
rect 252461 105571 252527 105574
rect 307477 105498 307543 105501
rect 307477 105496 310132 105498
rect 307477 105440 307482 105496
rect 307538 105440 310132 105496
rect 321510 105468 321570 105979
rect 307477 105438 310132 105440
rect 307477 105435 307543 105438
rect 305913 105226 305979 105229
rect 307661 105226 307727 105229
rect 305913 105224 307727 105226
rect 305913 105168 305918 105224
rect 305974 105168 307666 105224
rect 307722 105168 307727 105224
rect 305913 105166 307727 105168
rect 305913 105163 305979 105166
rect 307661 105163 307727 105166
rect 251725 105090 251791 105093
rect 248860 105088 251791 105090
rect 248860 105032 251730 105088
rect 251786 105032 251791 105088
rect 248860 105030 251791 105032
rect 251725 105027 251791 105030
rect 307661 105090 307727 105093
rect 307661 105088 310132 105090
rect 307661 105032 307666 105088
rect 307722 105032 310132 105088
rect 307661 105030 310132 105032
rect 307661 105027 307727 105030
rect 213913 104954 213979 104957
rect 213913 104952 217212 104954
rect 213913 104896 213918 104952
rect 213974 104896 217212 104952
rect 213913 104894 217212 104896
rect 213913 104891 213979 104894
rect 252185 104682 252251 104685
rect 248860 104680 252251 104682
rect 248860 104624 252190 104680
rect 252246 104624 252251 104680
rect 248860 104622 252251 104624
rect 252185 104619 252251 104622
rect 307569 104682 307635 104685
rect 307569 104680 310132 104682
rect 307569 104624 307574 104680
rect 307630 104624 310132 104680
rect 307569 104622 310132 104624
rect 307569 104619 307635 104622
rect 321694 104277 321754 104788
rect 214005 104274 214071 104277
rect 307477 104274 307543 104277
rect 214005 104272 217212 104274
rect 214005 104216 214010 104272
rect 214066 104216 217212 104272
rect 214005 104214 217212 104216
rect 307477 104272 310132 104274
rect 307477 104216 307482 104272
rect 307538 104216 310132 104272
rect 307477 104214 310132 104216
rect 321694 104272 321803 104277
rect 321694 104216 321742 104272
rect 321798 104216 321803 104272
rect 321694 104214 321803 104216
rect 214005 104211 214071 104214
rect 307477 104211 307543 104214
rect 321737 104211 321803 104214
rect 252369 104138 252435 104141
rect 248860 104136 252435 104138
rect 248860 104080 252374 104136
rect 252430 104080 252435 104136
rect 248860 104078 252435 104080
rect 252369 104075 252435 104078
rect 324313 104002 324379 104005
rect 321908 104000 324379 104002
rect 321908 103944 324318 104000
rect 324374 103944 324379 104000
rect 321908 103942 324379 103944
rect 324313 103939 324379 103942
rect 307661 103866 307727 103869
rect 307661 103864 310132 103866
rect 307661 103808 307666 103864
rect 307722 103808 310132 103864
rect 307661 103806 310132 103808
rect 307661 103803 307727 103806
rect 252461 103730 252527 103733
rect 248860 103728 252527 103730
rect 248860 103672 252466 103728
rect 252522 103672 252527 103728
rect 248860 103670 252527 103672
rect 252461 103667 252527 103670
rect 213913 103594 213979 103597
rect 213913 103592 217212 103594
rect 213913 103536 213918 103592
rect 213974 103536 217212 103592
rect 213913 103534 217212 103536
rect 213913 103531 213979 103534
rect 306741 103458 306807 103461
rect 306741 103456 310132 103458
rect 306741 103400 306746 103456
rect 306802 103400 310132 103456
rect 306741 103398 310132 103400
rect 306741 103395 306807 103398
rect 252277 103186 252343 103189
rect 324313 103186 324379 103189
rect 248860 103184 252343 103186
rect 248860 103128 252282 103184
rect 252338 103128 252343 103184
rect 248860 103126 252343 103128
rect 321908 103184 324379 103186
rect 321908 103128 324318 103184
rect 324374 103128 324379 103184
rect 321908 103126 324379 103128
rect 252277 103123 252343 103126
rect 324313 103123 324379 103126
rect 307477 103050 307543 103053
rect 307477 103048 310132 103050
rect 307477 102992 307482 103048
rect 307538 102992 310132 103048
rect 307477 102990 310132 102992
rect 307477 102987 307543 102990
rect 214741 102914 214807 102917
rect 214741 102912 217212 102914
rect 214741 102856 214746 102912
rect 214802 102856 217212 102912
rect 214741 102854 217212 102856
rect 214741 102851 214807 102854
rect 251173 102778 251239 102781
rect 248860 102776 251239 102778
rect 248860 102720 251178 102776
rect 251234 102720 251239 102776
rect 248860 102718 251239 102720
rect 251173 102715 251239 102718
rect 307661 102506 307727 102509
rect 307661 102504 310132 102506
rect 307661 102448 307666 102504
rect 307722 102448 310132 102504
rect 307661 102446 310132 102448
rect 307661 102443 307727 102446
rect 68142 102316 68816 102376
rect 64689 102234 64755 102237
rect 68142 102234 68202 102316
rect 64689 102232 68202 102234
rect 64689 102176 64694 102232
rect 64750 102176 68202 102232
rect 64689 102174 68202 102176
rect 64689 102171 64755 102174
rect 321510 102237 321570 102476
rect 213913 102234 213979 102237
rect 252461 102234 252527 102237
rect 213913 102232 217212 102234
rect 213913 102176 213918 102232
rect 213974 102176 217212 102232
rect 213913 102174 217212 102176
rect 248860 102232 252527 102234
rect 248860 102176 252466 102232
rect 252522 102176 252527 102232
rect 248860 102174 252527 102176
rect 321510 102232 321619 102237
rect 321510 102176 321558 102232
rect 321614 102176 321619 102232
rect 321510 102174 321619 102176
rect 213913 102171 213979 102174
rect 252461 102171 252527 102174
rect 321553 102171 321619 102174
rect 308213 102098 308279 102101
rect 308213 102096 310132 102098
rect 308213 102040 308218 102096
rect 308274 102040 310132 102096
rect 308213 102038 310132 102040
rect 308213 102035 308279 102038
rect 251909 101826 251975 101829
rect 248860 101824 251975 101826
rect 248860 101768 251914 101824
rect 251970 101768 251975 101824
rect 248860 101766 251975 101768
rect 251909 101763 251975 101766
rect 306557 101690 306623 101693
rect 324313 101690 324379 101693
rect 306557 101688 310132 101690
rect 306557 101632 306562 101688
rect 306618 101632 310132 101688
rect 306557 101630 310132 101632
rect 321908 101688 324379 101690
rect 321908 101632 324318 101688
rect 324374 101632 324379 101688
rect 321908 101630 324379 101632
rect 306557 101627 306623 101630
rect 324313 101627 324379 101630
rect 214925 101554 214991 101557
rect 214925 101552 217212 101554
rect 214925 101496 214930 101552
rect 214986 101496 217212 101552
rect 214925 101494 217212 101496
rect 214925 101491 214991 101494
rect 251173 101418 251239 101421
rect 248860 101416 251239 101418
rect 248860 101360 251178 101416
rect 251234 101360 251239 101416
rect 248860 101358 251239 101360
rect 251173 101355 251239 101358
rect 305678 101220 305684 101284
rect 305748 101282 305754 101284
rect 305748 101222 310132 101282
rect 305748 101220 305754 101222
rect 302734 101084 302740 101148
rect 302804 101146 302810 101148
rect 308213 101146 308279 101149
rect 302804 101144 308279 101146
rect 302804 101088 308218 101144
rect 308274 101088 308279 101144
rect 302804 101086 308279 101088
rect 302804 101084 302810 101086
rect 308213 101083 308279 101086
rect 213913 101010 213979 101013
rect 213913 101008 217212 101010
rect 213913 100952 213918 101008
rect 213974 100952 217212 101008
rect 213913 100950 217212 100952
rect 213913 100947 213979 100950
rect 252461 100874 252527 100877
rect 248860 100872 252527 100874
rect 248860 100816 252466 100872
rect 252522 100816 252527 100872
rect 248860 100814 252527 100816
rect 252461 100811 252527 100814
rect 307661 100874 307727 100877
rect 322933 100874 322999 100877
rect 307661 100872 310132 100874
rect 307661 100816 307666 100872
rect 307722 100816 310132 100872
rect 307661 100814 310132 100816
rect 321908 100872 322999 100874
rect 321908 100816 322938 100872
rect 322994 100816 322999 100872
rect 321908 100814 322999 100816
rect 307661 100811 307727 100814
rect 322933 100811 322999 100814
rect 67633 100738 67699 100741
rect 68142 100738 68816 100744
rect 67633 100736 68816 100738
rect 67633 100680 67638 100736
rect 67694 100684 68816 100736
rect 67694 100680 68202 100684
rect 67633 100678 68202 100680
rect 67633 100675 67699 100678
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 251541 100466 251607 100469
rect 248860 100464 251607 100466
rect 248860 100408 251546 100464
rect 251602 100408 251607 100464
rect 248860 100406 251607 100408
rect 251541 100403 251607 100406
rect 307569 100466 307635 100469
rect 307569 100464 310132 100466
rect 307569 100408 307574 100464
rect 307630 100408 310132 100464
rect 307569 100406 310132 100408
rect 307569 100403 307635 100406
rect 214005 100330 214071 100333
rect 214005 100328 217212 100330
rect 214005 100272 214010 100328
rect 214066 100272 217212 100328
rect 214005 100270 217212 100272
rect 214005 100267 214071 100270
rect 324497 100194 324563 100197
rect 321908 100192 324563 100194
rect 321908 100136 324502 100192
rect 324558 100136 324563 100192
rect 321908 100134 324563 100136
rect 324497 100131 324563 100134
rect 301630 99996 301636 100060
rect 301700 100058 301706 100060
rect 301700 99998 310132 100058
rect 301700 99996 301706 99998
rect 252001 99922 252067 99925
rect 248860 99920 252067 99922
rect 248860 99864 252006 99920
rect 252062 99864 252067 99920
rect 248860 99862 252067 99864
rect 252001 99859 252067 99862
rect 213913 99650 213979 99653
rect 307661 99650 307727 99653
rect 213913 99648 217212 99650
rect 213913 99592 213918 99648
rect 213974 99592 217212 99648
rect 213913 99590 217212 99592
rect 307661 99648 310132 99650
rect 307661 99592 307666 99648
rect 307722 99592 310132 99648
rect 307661 99590 310132 99592
rect 213913 99587 213979 99590
rect 307661 99587 307727 99590
rect 252461 99514 252527 99517
rect 248860 99512 252527 99514
rect 248860 99456 252466 99512
rect 252522 99456 252527 99512
rect 248860 99454 252527 99456
rect 252461 99451 252527 99454
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 324405 99378 324471 99381
rect 321908 99376 324471 99378
rect 321908 99320 324410 99376
rect 324466 99320 324471 99376
rect 583520 99364 584960 99454
rect 321908 99318 324471 99320
rect 324405 99315 324471 99318
rect 307661 99106 307727 99109
rect 307661 99104 310132 99106
rect 307661 99048 307666 99104
rect 307722 99048 310132 99104
rect 307661 99046 310132 99048
rect 307661 99043 307727 99046
rect 214005 98970 214071 98973
rect 251357 98970 251423 98973
rect 214005 98968 217212 98970
rect 214005 98912 214010 98968
rect 214066 98912 217212 98968
rect 214005 98910 217212 98912
rect 248860 98968 251423 98970
rect 248860 98912 251362 98968
rect 251418 98912 251423 98968
rect 248860 98910 251423 98912
rect 214005 98907 214071 98910
rect 251357 98907 251423 98910
rect 307569 98698 307635 98701
rect 307569 98696 310132 98698
rect 307569 98640 307574 98696
rect 307630 98640 310132 98696
rect 307569 98638 310132 98640
rect 307569 98635 307635 98638
rect 252461 98562 252527 98565
rect 248860 98560 252527 98562
rect 248860 98504 252466 98560
rect 252522 98504 252527 98560
rect 248860 98502 252527 98504
rect 252461 98499 252527 98502
rect 213913 98290 213979 98293
rect 307477 98290 307543 98293
rect 213913 98288 217212 98290
rect 213913 98232 213918 98288
rect 213974 98232 217212 98288
rect 213913 98230 217212 98232
rect 307477 98288 310132 98290
rect 307477 98232 307482 98288
rect 307538 98232 310132 98288
rect 307477 98230 310132 98232
rect 213913 98227 213979 98230
rect 307477 98227 307543 98230
rect 321878 98157 321938 98532
rect 321829 98152 321938 98157
rect 321829 98096 321834 98152
rect 321890 98096 321938 98152
rect 321829 98094 321938 98096
rect 321829 98091 321895 98094
rect 251950 98018 251956 98020
rect 248860 97958 251956 98018
rect 251950 97956 251956 97958
rect 252020 97956 252026 98020
rect 306741 97882 306807 97885
rect 306741 97880 310132 97882
rect 306741 97824 306746 97880
rect 306802 97824 310132 97880
rect 306741 97822 310132 97824
rect 306741 97819 306807 97822
rect 213913 97610 213979 97613
rect 261334 97610 261340 97612
rect 213913 97608 217212 97610
rect 213913 97552 213918 97608
rect 213974 97552 217212 97608
rect 213913 97550 217212 97552
rect 248860 97550 261340 97610
rect 213913 97547 213979 97550
rect 261334 97548 261340 97550
rect 261404 97548 261410 97612
rect 307477 97474 307543 97477
rect 307477 97472 310132 97474
rect 307477 97416 307482 97472
rect 307538 97416 310132 97472
rect 307477 97414 310132 97416
rect 307477 97411 307543 97414
rect 321369 97338 321435 97341
rect 321510 97338 321570 97852
rect 321369 97336 321570 97338
rect 321369 97280 321374 97336
rect 321430 97280 321570 97336
rect 321369 97278 321570 97280
rect 321369 97275 321435 97278
rect 166390 97140 166396 97204
rect 166460 97202 166466 97204
rect 214373 97202 214439 97205
rect 166460 97200 214439 97202
rect 166460 97144 214378 97200
rect 214434 97144 214439 97200
rect 166460 97142 214439 97144
rect 166460 97140 166466 97142
rect 214373 97139 214439 97142
rect 250110 97066 250116 97068
rect 248860 97006 250116 97066
rect 250110 97004 250116 97006
rect 250180 97066 250186 97068
rect 252185 97066 252251 97069
rect 250180 97064 252251 97066
rect 250180 97008 252190 97064
rect 252246 97008 252251 97064
rect 250180 97006 252251 97008
rect 250180 97004 250186 97006
rect 252185 97003 252251 97006
rect 306966 97004 306972 97068
rect 307036 97066 307042 97068
rect 324589 97066 324655 97069
rect 307036 97006 310132 97066
rect 321908 97064 324655 97066
rect 321908 97008 324594 97064
rect 324650 97008 324655 97064
rect 321908 97006 324655 97008
rect 307036 97004 307042 97006
rect 324589 97003 324655 97006
rect 214833 96930 214899 96933
rect 214833 96928 217212 96930
rect 214833 96872 214838 96928
rect 214894 96872 217212 96928
rect 214833 96870 217212 96872
rect 214833 96867 214899 96870
rect 251173 96658 251239 96661
rect 248860 96656 251239 96658
rect 248860 96600 251178 96656
rect 251234 96600 251239 96656
rect 248860 96598 251239 96600
rect 251173 96595 251239 96598
rect 307661 96658 307727 96661
rect 307661 96656 310132 96658
rect 307661 96600 307666 96656
rect 307722 96600 310132 96656
rect 307661 96598 310132 96600
rect 307661 96595 307727 96598
rect 214649 96386 214715 96389
rect 214649 96384 217212 96386
rect 214649 96328 214654 96384
rect 214710 96328 217212 96384
rect 214649 96326 217212 96328
rect 214649 96323 214715 96326
rect 251357 96250 251423 96253
rect 248860 96248 251423 96250
rect 248860 96192 251362 96248
rect 251418 96192 251423 96248
rect 248860 96190 251423 96192
rect 251357 96187 251423 96190
rect 307201 96250 307267 96253
rect 307201 96248 310132 96250
rect 307201 96192 307206 96248
rect 307262 96192 310132 96248
rect 307201 96190 310132 96192
rect 307201 96187 307267 96190
rect 171726 95916 171732 95980
rect 171796 95978 171802 95980
rect 321369 95978 321435 95981
rect 171796 95976 321435 95978
rect 171796 95920 321374 95976
rect 321430 95920 321435 95976
rect 171796 95918 321435 95920
rect 171796 95916 171802 95918
rect 321369 95915 321435 95918
rect 321510 95845 321570 96356
rect 321461 95840 321570 95845
rect 321461 95784 321466 95840
rect 321522 95784 321570 95840
rect 321461 95782 321570 95784
rect 321461 95779 321527 95782
rect 67541 94890 67607 94893
rect 194041 94890 194107 94893
rect 67541 94888 194107 94890
rect 67541 94832 67546 94888
rect 67602 94832 194046 94888
rect 194102 94832 194107 94888
rect 67541 94830 194107 94832
rect 67541 94827 67607 94830
rect 194041 94827 194107 94830
rect 109033 94756 109099 94757
rect 113725 94756 113791 94757
rect 131941 94756 132007 94757
rect 109033 94754 109062 94756
rect 108970 94752 109062 94754
rect 108970 94696 109038 94752
rect 108970 94694 109062 94696
rect 109033 94692 109062 94694
rect 109126 94692 109132 94756
rect 113680 94692 113686 94756
rect 113750 94754 113791 94756
rect 113750 94752 113842 94754
rect 113786 94696 113842 94752
rect 113750 94694 113842 94696
rect 113750 94692 113791 94694
rect 131904 94692 131910 94756
rect 131974 94754 132007 94756
rect 151721 94756 151787 94757
rect 151905 94756 151971 94757
rect 151721 94754 151766 94756
rect 131974 94752 132066 94754
rect 132002 94696 132066 94752
rect 131974 94694 132066 94696
rect 151674 94752 151766 94754
rect 151674 94696 151726 94752
rect 151674 94694 151766 94696
rect 131974 94692 132007 94694
rect 109033 94691 109099 94692
rect 113725 94691 113791 94692
rect 131941 94691 132007 94692
rect 151721 94692 151766 94694
rect 151830 94692 151836 94756
rect 151896 94692 151902 94756
rect 151966 94754 151972 94756
rect 151966 94694 152058 94754
rect 151966 94692 151972 94694
rect 151721 94691 151787 94692
rect 151905 94691 151971 94692
rect 114318 93876 114324 93940
rect 114388 93938 114394 93940
rect 172053 93938 172119 93941
rect 114388 93936 172119 93938
rect 114388 93880 172058 93936
rect 172114 93880 172119 93936
rect 114388 93878 172119 93880
rect 114388 93876 114394 93878
rect 172053 93875 172119 93878
rect 108062 93740 108068 93804
rect 108132 93802 108138 93804
rect 167678 93802 167684 93804
rect 108132 93742 167684 93802
rect 108132 93740 108138 93742
rect 167678 93740 167684 93742
rect 167748 93740 167754 93804
rect 173566 93740 173572 93804
rect 173636 93802 173642 93804
rect 324405 93802 324471 93805
rect 173636 93800 324471 93802
rect 173636 93744 324410 93800
rect 324466 93744 324471 93800
rect 173636 93742 324471 93744
rect 173636 93740 173642 93742
rect 324405 93739 324471 93742
rect 121729 93668 121795 93669
rect 121678 93666 121684 93668
rect 121638 93606 121684 93666
rect 121748 93664 121795 93668
rect 121790 93608 121795 93664
rect 121678 93604 121684 93606
rect 121748 93604 121795 93608
rect 121729 93603 121795 93604
rect 102041 93532 102107 93533
rect 107745 93532 107811 93533
rect 124489 93532 124555 93533
rect 101990 93530 101996 93532
rect 101950 93470 101996 93530
rect 102060 93528 102107 93532
rect 107694 93530 107700 93532
rect 102102 93472 102107 93528
rect 101990 93468 101996 93470
rect 102060 93468 102107 93472
rect 107654 93470 107700 93530
rect 107764 93528 107811 93532
rect 124438 93530 124444 93532
rect 107806 93472 107811 93528
rect 107694 93468 107700 93470
rect 107764 93468 107811 93472
rect 124398 93470 124444 93530
rect 124508 93528 124555 93532
rect 124550 93472 124555 93528
rect 124438 93468 124444 93470
rect 124508 93468 124555 93472
rect 102041 93467 102107 93468
rect 107745 93467 107811 93468
rect 124489 93467 124555 93468
rect 110137 93260 110203 93261
rect 119337 93260 119403 93261
rect 110086 93258 110092 93260
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 119286 93258 119292 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 119246 93198 119292 93258
rect 119356 93256 119403 93260
rect 119398 93200 119403 93256
rect 119286 93196 119292 93198
rect 119356 93196 119403 93200
rect 110137 93195 110203 93196
rect 119337 93195 119403 93196
rect 74809 92444 74875 92445
rect 74758 92442 74764 92444
rect 74718 92382 74764 92442
rect 74828 92440 74875 92444
rect 74870 92384 74875 92440
rect 74758 92380 74764 92382
rect 74828 92380 74875 92384
rect 85614 92380 85620 92444
rect 85684 92442 85690 92444
rect 85941 92442 86007 92445
rect 85684 92440 86007 92442
rect 85684 92384 85946 92440
rect 86002 92384 86007 92440
rect 85684 92382 86007 92384
rect 85684 92380 85690 92382
rect 74809 92379 74875 92380
rect 85941 92379 86007 92382
rect 93894 92380 93900 92444
rect 93964 92442 93970 92444
rect 94221 92442 94287 92445
rect 101857 92444 101923 92445
rect 101806 92442 101812 92444
rect 93964 92440 94287 92442
rect 93964 92384 94226 92440
rect 94282 92384 94287 92440
rect 93964 92382 94287 92384
rect 101766 92382 101812 92442
rect 101876 92440 101923 92444
rect 101918 92384 101923 92440
rect 93964 92380 93970 92382
rect 94221 92379 94287 92382
rect 101806 92380 101812 92382
rect 101876 92380 101923 92384
rect 115054 92380 115060 92444
rect 115124 92442 115130 92444
rect 115197 92442 115263 92445
rect 115473 92444 115539 92445
rect 115422 92442 115428 92444
rect 115124 92440 115263 92442
rect 115124 92384 115202 92440
rect 115258 92384 115263 92440
rect 115124 92382 115263 92384
rect 115382 92382 115428 92442
rect 115492 92440 115539 92444
rect 115534 92384 115539 92440
rect 115124 92380 115130 92382
rect 101857 92379 101923 92380
rect 115197 92379 115263 92382
rect 115422 92380 115428 92382
rect 115492 92380 115539 92384
rect 120206 92380 120212 92444
rect 120276 92442 120282 92444
rect 120349 92442 120415 92445
rect 124121 92444 124187 92445
rect 125961 92444 126027 92445
rect 133137 92444 133203 92445
rect 151721 92444 151787 92445
rect 124070 92442 124076 92444
rect 120276 92440 120415 92442
rect 120276 92384 120354 92440
rect 120410 92384 120415 92440
rect 120276 92382 120415 92384
rect 124030 92382 124076 92442
rect 124140 92440 124187 92444
rect 125910 92442 125916 92444
rect 124182 92384 124187 92440
rect 120276 92380 120282 92382
rect 115473 92379 115539 92380
rect 120349 92379 120415 92382
rect 124070 92380 124076 92382
rect 124140 92380 124187 92384
rect 125870 92382 125916 92442
rect 125980 92440 126027 92444
rect 133086 92442 133092 92444
rect 126022 92384 126027 92440
rect 125910 92380 125916 92382
rect 125980 92380 126027 92384
rect 133046 92382 133092 92442
rect 133156 92440 133203 92444
rect 133198 92384 133203 92440
rect 133086 92380 133092 92382
rect 133156 92380 133203 92384
rect 151670 92380 151676 92444
rect 151740 92442 151787 92444
rect 151740 92440 151832 92442
rect 151782 92384 151832 92440
rect 151740 92382 151832 92384
rect 151740 92380 151787 92382
rect 174486 92380 174492 92444
rect 174556 92442 174562 92444
rect 324589 92442 324655 92445
rect 174556 92440 324655 92442
rect 174556 92384 324594 92440
rect 324650 92384 324655 92440
rect 174556 92382 324655 92384
rect 174556 92380 174562 92382
rect 124121 92379 124187 92380
rect 125961 92379 126027 92380
rect 133137 92379 133203 92380
rect 151721 92379 151787 92380
rect 324589 92379 324655 92382
rect 111926 92244 111932 92308
rect 111996 92306 112002 92308
rect 166390 92306 166396 92308
rect 111996 92246 166396 92306
rect 111996 92244 112002 92246
rect 166390 92244 166396 92246
rect 166460 92244 166466 92308
rect 106038 92108 106044 92172
rect 106108 92170 106114 92172
rect 173341 92170 173407 92173
rect 106108 92168 173407 92170
rect 106108 92112 173346 92168
rect 173402 92112 173407 92168
rect 106108 92110 173407 92112
rect 106108 92108 106114 92110
rect 173341 92107 173407 92110
rect 88926 91700 88932 91764
rect 88996 91762 89002 91764
rect 89069 91762 89135 91765
rect 112345 91764 112411 91765
rect 112294 91762 112300 91764
rect 88996 91760 89135 91762
rect 88996 91704 89074 91760
rect 89130 91704 89135 91760
rect 88996 91702 89135 91704
rect 112254 91702 112300 91762
rect 112364 91760 112411 91764
rect 112406 91704 112411 91760
rect 88996 91700 89002 91702
rect 89069 91699 89135 91702
rect 112294 91700 112300 91702
rect 112364 91700 112411 91704
rect 122966 91700 122972 91764
rect 123036 91762 123042 91764
rect 123937 91762 124003 91765
rect 123036 91760 124003 91762
rect 123036 91704 123942 91760
rect 123998 91704 124003 91760
rect 123036 91702 124003 91704
rect 123036 91700 123042 91702
rect 112345 91699 112411 91700
rect 123937 91699 124003 91702
rect 151302 91700 151308 91764
rect 151372 91762 151378 91764
rect 151721 91762 151787 91765
rect 151372 91760 151787 91762
rect 151372 91704 151726 91760
rect 151782 91704 151787 91760
rect 151372 91702 151787 91704
rect 151372 91700 151378 91702
rect 151721 91699 151787 91702
rect 104198 91564 104204 91628
rect 104268 91626 104274 91628
rect 104525 91626 104591 91629
rect 104268 91624 104591 91626
rect 104268 91568 104530 91624
rect 104586 91568 104591 91624
rect 104268 91566 104591 91568
rect 104268 91564 104274 91566
rect 104525 91563 104591 91566
rect 106774 91564 106780 91628
rect 106844 91626 106850 91628
rect 106917 91626 106983 91629
rect 106844 91624 106983 91626
rect 106844 91568 106922 91624
rect 106978 91568 106983 91624
rect 106844 91566 106983 91568
rect 106844 91564 106850 91566
rect 106917 91563 106983 91566
rect 126462 91564 126468 91628
rect 126532 91626 126538 91628
rect 126605 91626 126671 91629
rect 126532 91624 126671 91626
rect 126532 91568 126610 91624
rect 126666 91568 126671 91624
rect 126532 91566 126671 91568
rect 126532 91564 126538 91566
rect 126605 91563 126671 91566
rect 98494 91428 98500 91492
rect 98564 91490 98570 91492
rect 99281 91490 99347 91493
rect 122833 91492 122899 91493
rect 98564 91488 99347 91490
rect 98564 91432 99286 91488
rect 99342 91432 99347 91488
rect 98564 91430 99347 91432
rect 98564 91428 98570 91430
rect 99281 91427 99347 91430
rect 122782 91428 122788 91492
rect 122852 91490 122899 91492
rect 122852 91488 122944 91490
rect 122894 91432 122944 91488
rect 122852 91430 122944 91432
rect 122852 91428 122899 91430
rect 122833 91427 122899 91428
rect 97022 91292 97028 91356
rect 97092 91354 97098 91356
rect 97901 91354 97967 91357
rect 97092 91352 97967 91354
rect 97092 91296 97906 91352
rect 97962 91296 97967 91352
rect 97092 91294 97967 91296
rect 97092 91292 97098 91294
rect 97901 91291 97967 91294
rect 98126 91292 98132 91356
rect 98196 91354 98202 91356
rect 99097 91354 99163 91357
rect 118233 91356 118299 91357
rect 118182 91354 118188 91356
rect 98196 91352 99163 91354
rect 98196 91296 99102 91352
rect 99158 91296 99163 91352
rect 98196 91294 99163 91296
rect 118142 91294 118188 91354
rect 118252 91352 118299 91356
rect 118294 91296 118299 91352
rect 98196 91292 98202 91294
rect 99097 91291 99163 91294
rect 118182 91292 118188 91294
rect 118252 91292 118299 91296
rect 118233 91291 118299 91292
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85021 91218 85087 91221
rect 86769 91220 86835 91221
rect 86718 91218 86724 91220
rect 84396 91216 85087 91218
rect 84396 91160 85026 91216
rect 85082 91160 85087 91216
rect 84396 91158 85087 91160
rect 86678 91158 86724 91218
rect 86788 91216 86835 91220
rect 86830 91160 86835 91216
rect 84396 91156 84402 91158
rect 85021 91155 85087 91158
rect 86718 91156 86724 91158
rect 86788 91156 86835 91160
rect 87086 91156 87092 91220
rect 87156 91218 87162 91220
rect 87413 91218 87479 91221
rect 87156 91216 87479 91218
rect 87156 91160 87418 91216
rect 87474 91160 87479 91216
rect 87156 91158 87479 91160
rect 87156 91156 87162 91158
rect 86769 91155 86835 91156
rect 87413 91155 87479 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 91001 91218 91067 91221
rect 90284 91216 91067 91218
rect 90284 91160 91006 91216
rect 91062 91160 91067 91216
rect 90284 91158 91067 91160
rect 90284 91156 90290 91158
rect 91001 91155 91067 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92381 91218 92447 91221
rect 91388 91216 92447 91218
rect 91388 91160 92386 91216
rect 92442 91160 92447 91216
rect 91388 91158 92447 91160
rect 91388 91156 91394 91158
rect 92381 91155 92447 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 95049 91220 95115 91221
rect 94998 91218 95004 91220
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 94958 91158 95004 91218
rect 95068 91216 95115 91220
rect 95110 91160 95115 91216
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 94998 91156 95004 91158
rect 95068 91156 95115 91160
rect 96102 91156 96108 91220
rect 96172 91218 96178 91220
rect 96521 91218 96587 91221
rect 96172 91216 96587 91218
rect 96172 91160 96526 91216
rect 96582 91160 96587 91216
rect 96172 91158 96587 91160
rect 96172 91156 96178 91158
rect 95049 91155 95115 91156
rect 96521 91155 96587 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97809 91218 97875 91221
rect 99189 91220 99255 91221
rect 99189 91218 99236 91220
rect 97276 91216 97875 91218
rect 97276 91160 97814 91216
rect 97870 91160 97875 91216
rect 97276 91158 97875 91160
rect 99144 91216 99236 91218
rect 99144 91160 99194 91216
rect 99144 91158 99236 91160
rect 97276 91156 97282 91158
rect 97809 91155 97875 91158
rect 99189 91156 99236 91158
rect 99300 91156 99306 91220
rect 99598 91156 99604 91220
rect 99668 91218 99674 91220
rect 99925 91218 99991 91221
rect 99668 91216 99991 91218
rect 99668 91160 99930 91216
rect 99986 91160 99991 91216
rect 99668 91158 99991 91160
rect 99668 91156 99674 91158
rect 99189 91155 99255 91156
rect 99925 91155 99991 91158
rect 100518 91156 100524 91220
rect 100588 91218 100594 91220
rect 100661 91218 100727 91221
rect 100588 91216 100727 91218
rect 100588 91160 100666 91216
rect 100722 91160 100727 91216
rect 100588 91158 100727 91160
rect 100588 91156 100594 91158
rect 100661 91155 100727 91158
rect 101622 91156 101628 91220
rect 101692 91218 101698 91220
rect 102041 91218 102107 91221
rect 102961 91220 103027 91221
rect 102910 91218 102916 91220
rect 101692 91216 102107 91218
rect 101692 91160 102046 91216
rect 102102 91160 102107 91216
rect 101692 91158 102107 91160
rect 102870 91158 102916 91218
rect 102980 91216 103027 91220
rect 103022 91160 103027 91216
rect 101692 91156 101698 91158
rect 102041 91155 102107 91158
rect 102910 91156 102916 91158
rect 102980 91156 103027 91160
rect 103278 91156 103284 91220
rect 103348 91218 103354 91220
rect 103421 91218 103487 91221
rect 104617 91220 104683 91221
rect 104566 91218 104572 91220
rect 103348 91216 103487 91218
rect 103348 91160 103426 91216
rect 103482 91160 103487 91216
rect 103348 91158 103487 91160
rect 104526 91158 104572 91218
rect 104636 91216 104683 91220
rect 104678 91160 104683 91216
rect 103348 91156 103354 91158
rect 102961 91155 103027 91156
rect 103421 91155 103487 91158
rect 104566 91156 104572 91158
rect 104636 91156 104683 91160
rect 105118 91156 105124 91220
rect 105188 91218 105194 91220
rect 106181 91218 106247 91221
rect 105188 91216 106247 91218
rect 105188 91160 106186 91216
rect 106242 91160 106247 91216
rect 105188 91158 106247 91160
rect 105188 91156 105194 91158
rect 104617 91155 104683 91156
rect 106181 91155 106247 91158
rect 106406 91156 106412 91220
rect 106476 91218 106482 91220
rect 106641 91218 106707 91221
rect 106476 91216 106707 91218
rect 106476 91160 106646 91216
rect 106702 91160 106707 91216
rect 106476 91158 106707 91160
rect 106476 91156 106482 91158
rect 106641 91155 106707 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110321 91218 110387 91221
rect 110689 91220 110755 91221
rect 110638 91218 110644 91220
rect 109604 91216 110387 91218
rect 109604 91160 110326 91216
rect 110382 91160 110387 91216
rect 109604 91158 110387 91160
rect 110598 91158 110644 91218
rect 110708 91216 110755 91220
rect 110750 91160 110755 91216
rect 109604 91156 109610 91158
rect 110321 91155 110387 91158
rect 110638 91156 110644 91158
rect 110708 91156 110755 91160
rect 111190 91156 111196 91220
rect 111260 91218 111266 91220
rect 111701 91218 111767 91221
rect 111260 91216 111767 91218
rect 111260 91160 111706 91216
rect 111762 91160 111767 91216
rect 111260 91158 111767 91160
rect 111260 91156 111266 91158
rect 110689 91155 110755 91156
rect 111701 91155 111767 91158
rect 113214 91156 113220 91220
rect 113284 91218 113290 91220
rect 114461 91218 114527 91221
rect 115749 91220 115815 91221
rect 116761 91220 116827 91221
rect 117129 91220 117195 91221
rect 115749 91218 115796 91220
rect 113284 91216 114527 91218
rect 113284 91160 114466 91216
rect 114522 91160 114527 91216
rect 113284 91158 114527 91160
rect 115704 91216 115796 91218
rect 115704 91160 115754 91216
rect 115704 91158 115796 91160
rect 113284 91156 113290 91158
rect 114461 91155 114527 91158
rect 115749 91156 115796 91158
rect 115860 91156 115866 91220
rect 116710 91218 116716 91220
rect 116670 91158 116716 91218
rect 116780 91216 116827 91220
rect 117078 91218 117084 91220
rect 116822 91160 116827 91216
rect 116710 91156 116716 91158
rect 116780 91156 116827 91160
rect 117038 91158 117084 91218
rect 117148 91216 117195 91220
rect 117190 91160 117195 91216
rect 117078 91156 117084 91158
rect 117148 91156 117195 91160
rect 117998 91156 118004 91220
rect 118068 91218 118074 91220
rect 118601 91218 118667 91221
rect 118068 91216 118667 91218
rect 118068 91160 118606 91216
rect 118662 91160 118667 91216
rect 118068 91158 118667 91160
rect 118068 91156 118074 91158
rect 115749 91155 115815 91156
rect 116761 91155 116827 91156
rect 117129 91155 117195 91156
rect 118601 91155 118667 91158
rect 119654 91156 119660 91220
rect 119724 91218 119730 91220
rect 119981 91218 120047 91221
rect 119724 91216 120047 91218
rect 119724 91160 119986 91216
rect 120042 91160 120047 91216
rect 119724 91158 120047 91160
rect 119724 91156 119730 91158
rect 119981 91155 120047 91158
rect 120574 91156 120580 91220
rect 120644 91218 120650 91220
rect 121085 91218 121151 91221
rect 120644 91216 121151 91218
rect 120644 91160 121090 91216
rect 121146 91160 121151 91216
rect 120644 91158 121151 91160
rect 120644 91156 120650 91158
rect 121085 91155 121151 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122373 91218 122439 91221
rect 122116 91216 122439 91218
rect 122116 91160 122378 91216
rect 122434 91160 122439 91216
rect 122116 91158 122439 91160
rect 122116 91156 122122 91158
rect 122373 91155 122439 91158
rect 125358 91156 125364 91220
rect 125428 91218 125434 91220
rect 125501 91218 125567 91221
rect 125428 91216 125567 91218
rect 125428 91160 125506 91216
rect 125562 91160 125567 91216
rect 125428 91158 125567 91160
rect 125428 91156 125434 91158
rect 125501 91155 125567 91158
rect 126646 91156 126652 91220
rect 126716 91218 126722 91220
rect 126881 91218 126947 91221
rect 126716 91216 126947 91218
rect 126716 91160 126886 91216
rect 126942 91160 126947 91216
rect 126716 91158 126947 91160
rect 126716 91156 126722 91158
rect 126881 91155 126947 91158
rect 127566 91156 127572 91220
rect 127636 91156 127642 91220
rect 129406 91156 129412 91220
rect 129476 91218 129482 91220
rect 129641 91218 129707 91221
rect 129476 91216 129707 91218
rect 129476 91160 129646 91216
rect 129702 91160 129707 91216
rect 129476 91158 129707 91160
rect 129476 91156 129482 91158
rect 127574 91082 127634 91156
rect 129641 91155 129707 91158
rect 130694 91156 130700 91220
rect 130764 91218 130770 91220
rect 131021 91218 131087 91221
rect 130764 91216 131087 91218
rect 130764 91160 131026 91216
rect 131082 91160 131087 91216
rect 130764 91158 131087 91160
rect 130764 91156 130770 91158
rect 131021 91155 131087 91158
rect 134374 91156 134380 91220
rect 134444 91218 134450 91220
rect 135069 91218 135135 91221
rect 134444 91216 135135 91218
rect 134444 91160 135074 91216
rect 135130 91160 135135 91216
rect 134444 91158 135135 91160
rect 134444 91156 134450 91158
rect 135069 91155 135135 91158
rect 135662 91156 135668 91220
rect 135732 91218 135738 91220
rect 135897 91218 135963 91221
rect 135732 91216 135963 91218
rect 135732 91160 135902 91216
rect 135958 91160 135963 91216
rect 135732 91158 135963 91160
rect 135732 91156 135738 91158
rect 135897 91155 135963 91158
rect 167494 91082 167500 91084
rect 127574 91022 167500 91082
rect 167494 91020 167500 91022
rect 167564 91020 167570 91084
rect 67449 89722 67515 89725
rect 214741 89722 214807 89725
rect 67449 89720 214807 89722
rect 67449 89664 67454 89720
rect 67510 89664 214746 89720
rect 214802 89664 214807 89720
rect 67449 89662 214807 89664
rect 67449 89659 67515 89662
rect 214741 89659 214807 89662
rect 214557 89178 214623 89181
rect 307150 89178 307156 89180
rect 214557 89176 307156 89178
rect 214557 89120 214562 89176
rect 214618 89120 307156 89176
rect 214557 89118 307156 89120
rect 214557 89115 214623 89118
rect 307150 89116 307156 89118
rect 307220 89116 307226 89180
rect 178902 88980 178908 89044
rect 178972 89042 178978 89044
rect 331305 89042 331371 89045
rect 178972 89040 331371 89042
rect 178972 88984 331310 89040
rect 331366 88984 331371 89040
rect 178972 88982 331371 88984
rect 178972 88980 178978 88982
rect 331305 88979 331371 88982
rect 110689 88226 110755 88229
rect 166257 88226 166323 88229
rect 110689 88224 166323 88226
rect 110689 88168 110694 88224
rect 110750 88168 166262 88224
rect 166318 88168 166323 88224
rect 110689 88166 166323 88168
rect 110689 88163 110755 88166
rect 166257 88163 166323 88166
rect 104617 86866 104683 86869
rect 166206 86866 166212 86868
rect 104617 86864 166212 86866
rect 104617 86808 104622 86864
rect 104678 86808 166212 86864
rect 104617 86806 166212 86808
rect 104617 86803 104683 86806
rect 166206 86804 166212 86806
rect 166276 86804 166282 86868
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 110321 84146 110387 84149
rect 170254 84146 170260 84148
rect 110321 84144 170260 84146
rect 110321 84088 110326 84144
rect 110382 84088 170260 84144
rect 110321 84086 170260 84088
rect 110321 84083 110387 84086
rect 170254 84084 170260 84086
rect 170324 84084 170330 84148
rect 179638 79324 179644 79388
rect 179708 79386 179714 79388
rect 310513 79386 310579 79389
rect 179708 79384 310579 79386
rect 179708 79328 310518 79384
rect 310574 79328 310579 79384
rect 179708 79326 310579 79328
rect 179708 79324 179714 79326
rect 310513 79323 310579 79326
rect 99189 78570 99255 78573
rect 169150 78570 169156 78572
rect 99189 78568 169156 78570
rect 99189 78512 99194 78568
rect 99250 78512 169156 78568
rect 99189 78510 169156 78512
rect 99189 78507 99255 78510
rect 169150 78508 169156 78510
rect 169220 78508 169226 78572
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 88333 69594 88399 69597
rect 300158 69594 300164 69596
rect 88333 69592 300164 69594
rect 88333 69536 88338 69592
rect 88394 69536 300164 69592
rect 88333 69534 300164 69536
rect 88333 69531 88399 69534
rect 300158 69532 300164 69534
rect 300228 69532 300234 69596
rect 16573 62794 16639 62797
rect 301630 62794 301636 62796
rect 16573 62792 301636 62794
rect 16573 62736 16578 62792
rect 16634 62736 301636 62792
rect 16573 62734 301636 62736
rect 16573 62731 16639 62734
rect 301630 62732 301636 62734
rect 301700 62732 301706 62796
rect 13813 59938 13879 59941
rect 293166 59938 293172 59940
rect 13813 59936 293172 59938
rect 13813 59880 13818 59936
rect 13874 59880 293172 59936
rect 13813 59878 293172 59880
rect 13813 59875 13879 59878
rect 293166 59876 293172 59878
rect 293236 59876 293242 59940
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 52453 58578 52519 58581
rect 291694 58578 291700 58580
rect 52453 58576 291700 58578
rect 52453 58520 52458 58576
rect 52514 58520 291700 58576
rect 52453 58518 291700 58520
rect 52453 58515 52519 58518
rect 291694 58516 291700 58518
rect 291764 58516 291770 58580
rect 177062 50220 177068 50284
rect 177132 50282 177138 50284
rect 347773 50282 347839 50285
rect 177132 50280 347839 50282
rect 177132 50224 347778 50280
rect 347834 50224 347839 50280
rect 177132 50222 347839 50224
rect 177132 50220 177138 50222
rect 347773 50219 347839 50222
rect 35893 48922 35959 48925
rect 302734 48922 302740 48924
rect 35893 48920 302740 48922
rect 35893 48864 35898 48920
rect 35954 48864 302740 48920
rect 35893 48862 302740 48864
rect 35893 48859 35959 48862
rect 302734 48860 302740 48862
rect 302804 48860 302810 48924
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 176326 39204 176332 39268
rect 176396 39266 176402 39268
rect 579613 39266 579679 39269
rect 176396 39264 579679 39266
rect 176396 39208 579618 39264
rect 579674 39208 579679 39264
rect 176396 39206 579679 39208
rect 176396 39204 176402 39206
rect 579613 39203 579679 39206
rect 2773 37906 2839 37909
rect 305494 37906 305500 37908
rect 2773 37904 305500 37906
rect 2773 37848 2778 37904
rect 2834 37848 305500 37904
rect 2773 37846 305500 37848
rect 2773 37843 2839 37846
rect 305494 37844 305500 37846
rect 305564 37844 305570 37908
rect 579889 33146 579955 33149
rect 583520 33146 584960 33236
rect 579889 33144 584960 33146
rect 579889 33088 579894 33144
rect 579950 33088 584960 33144
rect 579889 33086 584960 33088
rect 579889 33083 579955 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 52545 26890 52611 26893
rect 295926 26890 295932 26892
rect 52545 26888 295932 26890
rect 52545 26832 52550 26888
rect 52606 26832 295932 26888
rect 52545 26830 295932 26832
rect 52545 26827 52611 26830
rect 295926 26828 295932 26830
rect 295996 26828 296002 26892
rect 179270 21252 179276 21316
rect 179340 21314 179346 21316
rect 332685 21314 332751 21317
rect 179340 21312 332751 21314
rect 179340 21256 332690 21312
rect 332746 21256 332751 21312
rect 179340 21254 332751 21256
rect 179340 21252 179346 21254
rect 332685 21251 332751 21254
rect 579889 19818 579955 19821
rect 583520 19818 584960 19908
rect 579889 19816 584960 19818
rect 579889 19760 579894 19816
rect 579950 19760 584960 19816
rect 579889 19758 584960 19760
rect 579889 19755 579955 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 184790 18668 184796 18732
rect 184860 18730 184866 18732
rect 345657 18730 345723 18733
rect 184860 18728 345723 18730
rect 184860 18672 345662 18728
rect 345718 18672 345723 18728
rect 184860 18670 345723 18672
rect 184860 18668 184866 18670
rect 345657 18667 345723 18670
rect 27613 18594 27679 18597
rect 275134 18594 275140 18596
rect 27613 18592 275140 18594
rect 27613 18536 27618 18592
rect 27674 18536 275140 18592
rect 27613 18534 275140 18536
rect 27613 18531 27679 18534
rect 275134 18532 275140 18534
rect 275204 18532 275210 18596
rect 2681 16554 2747 16557
rect 250110 16554 250116 16556
rect 2681 16552 250116 16554
rect 2681 16496 2686 16552
rect 2742 16496 250116 16552
rect 2681 16494 250116 16496
rect 2681 16491 2747 16494
rect 250110 16492 250116 16494
rect 250180 16492 250186 16556
rect 1393 15330 1459 15333
rect 2681 15330 2747 15333
rect 1393 15328 2747 15330
rect 1393 15272 1398 15328
rect 1454 15272 2686 15328
rect 2742 15272 2747 15328
rect 1393 15270 2747 15272
rect 1393 15267 1459 15270
rect 2681 15267 2747 15270
rect 30097 13018 30163 13021
rect 305678 13018 305684 13020
rect 30097 13016 305684 13018
rect 30097 12960 30102 13016
rect 30158 12960 305684 13016
rect 30097 12958 305684 12960
rect 30097 12955 30163 12958
rect 305678 12956 305684 12958
rect 305748 12956 305754 13020
rect 56593 8938 56659 8941
rect 306966 8938 306972 8940
rect 56593 8936 306972 8938
rect 56593 8880 56598 8936
rect 56654 8880 306972 8936
rect 56593 8878 306972 8880
rect 56593 8875 56659 8878
rect 306966 8876 306972 8878
rect 307036 8876 307042 8940
rect 582465 6626 582531 6629
rect 583520 6626 584960 6716
rect 582465 6624 584960 6626
rect -960 6490 480 6580
rect 582465 6568 582470 6624
rect 582526 6568 584960 6624
rect 582465 6566 584960 6568
rect 582465 6563 582531 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 175038 6156 175044 6220
rect 175108 6218 175114 6220
rect 301957 6218 302023 6221
rect 175108 6216 302023 6218
rect 175108 6160 301962 6216
rect 302018 6160 302023 6216
rect 175108 6158 302023 6160
rect 175108 6156 175114 6158
rect 301957 6155 302023 6158
rect 271086 3980 271092 4044
rect 271156 4042 271162 4044
rect 278313 4042 278379 4045
rect 271156 4040 278379 4042
rect 271156 3984 278318 4040
rect 278374 3984 278379 4040
rect 271156 3982 278379 3984
rect 271156 3980 271162 3982
rect 278313 3979 278379 3982
rect 296069 4042 296135 4045
rect 296478 4042 296484 4044
rect 296069 4040 296484 4042
rect 296069 3984 296074 4040
rect 296130 3984 296484 4040
rect 296069 3982 296484 3984
rect 296069 3979 296135 3982
rect 296478 3980 296484 3982
rect 296548 3980 296554 4044
rect 304206 3980 304212 4044
rect 304276 4042 304282 4044
rect 309041 4042 309107 4045
rect 304276 4040 309107 4042
rect 304276 3984 309046 4040
rect 309102 3984 309107 4040
rect 304276 3982 309107 3984
rect 304276 3980 304282 3982
rect 309041 3979 309107 3982
rect 301446 3572 301452 3636
rect 301516 3634 301522 3636
rect 319713 3634 319779 3637
rect 301516 3632 319779 3634
rect 301516 3576 319718 3632
rect 319774 3576 319779 3632
rect 301516 3574 319779 3576
rect 301516 3572 301522 3574
rect 319713 3571 319779 3574
rect 299974 3436 299980 3500
rect 300044 3498 300050 3500
rect 303153 3498 303219 3501
rect 300044 3496 303219 3498
rect 300044 3440 303158 3496
rect 303214 3440 303219 3496
rect 300044 3438 303219 3440
rect 300044 3436 300050 3438
rect 303153 3435 303219 3438
rect 307937 3498 308003 3501
rect 332542 3498 332548 3500
rect 307937 3496 332548 3498
rect 307937 3440 307942 3496
rect 307998 3440 332548 3496
rect 307937 3438 332548 3440
rect 307937 3435 308003 3438
rect 332542 3436 332548 3438
rect 332612 3436 332618 3500
rect 340822 3436 340828 3500
rect 340892 3498 340898 3500
rect 342161 3498 342227 3501
rect 340892 3496 342227 3498
rect 340892 3440 342166 3496
rect 342222 3440 342227 3496
rect 340892 3438 342227 3440
rect 340892 3436 340898 3438
rect 342161 3435 342227 3438
rect 125869 3362 125935 3365
rect 169702 3362 169708 3364
rect 125869 3360 169708 3362
rect 125869 3304 125874 3360
rect 125930 3304 169708 3360
rect 125869 3302 169708 3304
rect 125869 3299 125935 3302
rect 169702 3300 169708 3302
rect 169772 3300 169778 3364
rect 269614 3300 269620 3364
rect 269684 3362 269690 3364
rect 310237 3362 310303 3365
rect 269684 3360 310303 3362
rect 269684 3304 310242 3360
rect 310298 3304 310303 3360
rect 269684 3302 310303 3304
rect 269684 3300 269690 3302
rect 310237 3299 310303 3302
rect 176510 1940 176516 2004
rect 176580 2002 176586 2004
rect 339861 2002 339927 2005
rect 176580 2000 339927 2002
rect 176580 1944 339866 2000
rect 339922 1944 339927 2000
rect 176580 1942 339927 1944
rect 176580 1940 176586 1942
rect 339861 1939 339927 1942
<< obsm3 >>
rect 68800 171594 164756 174600
rect 68800 171534 164694 171594
rect 68800 129304 164756 171534
rect 68816 129244 164756 129304
rect 68800 128080 164756 129244
rect 68816 128020 164756 128080
rect 68800 126312 164756 128020
rect 68816 126252 164756 126312
rect 68800 125224 164756 126252
rect 68816 125164 164756 125224
rect 68800 123592 164756 125164
rect 68816 123532 164756 123592
rect 68800 122640 164756 123532
rect 68816 122580 164756 122640
rect 68800 120872 164756 122580
rect 68816 120812 164756 120872
rect 68800 111754 164756 120812
rect 68800 111694 164694 111754
rect 68800 110122 164756 111694
rect 68800 110062 164694 110122
rect 68800 108762 164756 110062
rect 68800 108702 164694 108762
rect 68800 102376 164756 108702
rect 68816 102316 164756 102376
rect 68800 100744 164756 102316
rect 68816 100684 164756 100744
rect 68800 95100 164756 100684
<< via3 >>
rect 243492 586468 243556 586532
rect 247172 585380 247236 585444
rect 243676 585168 243740 585172
rect 243676 585112 243690 585168
rect 243690 585112 243740 585168
rect 243676 585108 243740 585112
rect 63540 584564 63604 584628
rect 50844 583884 50908 583948
rect 58940 582524 59004 582588
rect 243676 580892 243740 580956
rect 243308 579532 243372 579596
rect 57836 579124 57900 579188
rect 243492 578852 243556 578916
rect 295380 578852 295444 578916
rect 60044 575724 60108 575788
rect 61884 572324 61948 572388
rect 246988 569604 247052 569668
rect 63540 558180 63604 558244
rect 54340 557500 54404 557564
rect 244228 553284 244292 553348
rect 244412 546484 244476 546548
rect 55628 532204 55692 532268
rect 245700 529484 245764 529548
rect 59124 525404 59188 525468
rect 63540 511804 63604 511868
rect 62068 510444 62132 510508
rect 245884 489364 245948 489428
rect 62068 485828 62132 485892
rect 63724 473180 63788 473244
rect 49556 469780 49620 469844
rect 328500 467876 328564 467940
rect 53604 464884 53668 464948
rect 331260 452644 331324 452708
rect 63724 449924 63788 449988
rect 63356 448564 63420 448628
rect 57652 434556 57716 434620
rect 53420 430612 53484 430676
rect 64092 429252 64156 429316
rect 63172 421364 63236 421428
rect 243308 407220 243372 407284
rect 53420 405588 53484 405652
rect 247172 405452 247236 405516
rect 57652 404908 57716 404972
rect 63172 404500 63236 404564
rect 61884 404364 61948 404428
rect 66852 403684 66916 403748
rect 243308 403548 243372 403612
rect 52500 401644 52564 401708
rect 245884 400964 245948 401028
rect 244412 400828 244476 400892
rect 58940 399468 59004 399532
rect 50844 398108 50908 398172
rect 63540 397972 63604 398036
rect 180012 389948 180076 390012
rect 244228 389812 244292 389876
rect 60044 386956 60108 387020
rect 178540 386956 178604 387020
rect 246988 380292 247052 380356
rect 242940 380156 243004 380220
rect 70900 378116 70964 378180
rect 295012 375260 295076 375324
rect 146892 368460 146956 368524
rect 295564 367644 295628 367708
rect 134380 367100 134444 367164
rect 332548 365740 332612 365804
rect 245700 362204 245764 362268
rect 340828 360164 340892 360228
rect 119660 359348 119724 359412
rect 172284 359348 172348 359412
rect 299980 358940 300044 359004
rect 296484 358804 296548 358868
rect 129044 357580 129108 357644
rect 298508 357580 298572 357644
rect 293908 357368 293972 357372
rect 293908 357312 293958 357368
rect 293958 357312 293972 357368
rect 293908 357308 293972 357312
rect 64092 356628 64156 356692
rect 301452 356356 301516 356420
rect 304212 356220 304276 356284
rect 292620 356084 292684 356148
rect 177068 355268 177132 355332
rect 53604 354588 53668 354652
rect 152412 352548 152476 352612
rect 179828 352548 179892 352612
rect 176516 350100 176580 350164
rect 178540 349692 178604 349756
rect 125732 341396 125796 341460
rect 176332 339220 176396 339284
rect 59124 327660 59188 327724
rect 179276 327660 179340 327724
rect 175044 321540 175108 321604
rect 49556 314740 49620 314804
rect 161980 314740 162044 314804
rect 295380 312156 295444 312220
rect 293172 309028 293236 309092
rect 293908 305356 293972 305420
rect 128860 304948 128924 305012
rect 148180 303588 148244 303652
rect 292620 303452 292684 303516
rect 124260 301412 124324 301476
rect 144684 301412 144748 301476
rect 152412 301140 152476 301204
rect 138612 301004 138676 301068
rect 130332 299508 130396 299572
rect 69060 298692 69124 298756
rect 153700 296924 153764 296988
rect 169708 295564 169772 295628
rect 160692 295428 160756 295492
rect 64644 294536 64708 294540
rect 64644 294480 64694 294536
rect 64694 294480 64708 294536
rect 64644 294476 64708 294480
rect 173572 294476 173636 294540
rect 174492 293932 174556 293996
rect 122052 292572 122116 292636
rect 120028 291892 120092 291956
rect 124076 290396 124140 290460
rect 129044 289172 129108 289236
rect 70532 288084 70596 288148
rect 124260 286996 124324 287060
rect 124260 286588 124324 286652
rect 120580 285908 120644 285972
rect 125732 285636 125796 285700
rect 54340 284276 54404 284340
rect 119660 283324 119724 283388
rect 126100 283188 126164 283252
rect 292620 281692 292684 281756
rect 179092 279516 179156 279580
rect 166396 275980 166460 276044
rect 149652 272580 149716 272644
rect 55628 271764 55692 271828
rect 171732 265508 171796 265572
rect 149652 264964 149716 265028
rect 177068 262108 177132 262172
rect 177068 259660 177132 259724
rect 64460 256804 64524 256868
rect 295380 257076 295444 257140
rect 179276 256668 179340 256732
rect 122052 255852 122116 255916
rect 149652 255852 149716 255916
rect 172284 255232 172348 255236
rect 172284 255176 172334 255232
rect 172334 255176 172348 255232
rect 172284 255172 172348 255176
rect 63172 254008 63236 254012
rect 63172 253952 63186 254008
rect 63186 253952 63236 254008
rect 63172 253948 63236 253952
rect 66852 252996 66916 253060
rect 67404 252996 67468 253060
rect 63356 252512 63420 252516
rect 63356 252456 63406 252512
rect 63406 252456 63420 252512
rect 63356 252452 63420 252456
rect 69060 252316 69124 252380
rect 295012 248236 295076 248300
rect 179276 248100 179340 248164
rect 295564 246256 295628 246260
rect 295564 246200 295578 246256
rect 295578 246200 295628 246256
rect 295564 246196 295628 246200
rect 61884 244428 61948 244492
rect 179644 243612 179708 243676
rect 144684 243476 144748 243540
rect 166212 243476 166276 243540
rect 179828 243476 179892 243540
rect 146892 242932 146956 242996
rect 152412 241708 152476 241772
rect 126100 241436 126164 241500
rect 298508 240756 298572 240820
rect 295380 240076 295444 240140
rect 292620 239184 292684 239188
rect 292620 239128 292670 239184
rect 292670 239128 292684 239184
rect 292620 239124 292684 239128
rect 124076 238716 124140 238780
rect 57836 238580 57900 238644
rect 161980 238580 162044 238644
rect 184796 237356 184860 237420
rect 61884 237220 61948 237284
rect 120580 237084 120644 237148
rect 134380 236948 134444 237012
rect 293172 235316 293236 235380
rect 64460 235180 64524 235244
rect 169708 231780 169772 231844
rect 179828 231840 179892 231844
rect 179828 231784 179842 231840
rect 179842 231784 179892 231840
rect 179828 231780 179892 231784
rect 331260 228924 331324 228988
rect 328684 227700 328748 227764
rect 179092 226884 179156 226948
rect 178908 226340 178972 226404
rect 256740 225524 256804 225588
rect 259500 224164 259564 224228
rect 338252 223620 338316 223684
rect 252508 222804 252572 222868
rect 63172 222124 63236 222188
rect 149652 221988 149716 222052
rect 166396 220764 166460 220828
rect 329788 220824 329852 220828
rect 329788 220768 329838 220824
rect 329838 220768 329852 220824
rect 329788 220764 329852 220768
rect 327028 219328 327092 219332
rect 327028 219272 327078 219328
rect 327078 219272 327092 219328
rect 327028 219268 327092 219272
rect 130332 213148 130396 213212
rect 336780 213148 336844 213212
rect 119844 210292 119908 210356
rect 265020 204852 265084 204916
rect 260972 202268 261036 202332
rect 128860 202132 128924 202196
rect 266308 200772 266372 200836
rect 64644 200636 64708 200700
rect 327580 196692 327644 196756
rect 138612 196556 138676 196620
rect 345060 196556 345124 196620
rect 335676 195196 335740 195260
rect 257844 193972 257908 194036
rect 67404 193836 67468 193900
rect 263732 192476 263796 192540
rect 269620 191116 269684 191180
rect 260788 190980 260852 191044
rect 271092 188532 271156 188596
rect 263548 188396 263612 188460
rect 148180 188260 148244 188324
rect 318012 186900 318076 186964
rect 255452 186356 255516 186420
rect 320220 185540 320284 185604
rect 153700 184180 153764 184244
rect 265204 182820 265268 182884
rect 166396 182140 166460 182204
rect 169708 181596 169772 181660
rect 255268 181460 255332 181524
rect 322060 181324 322124 181388
rect 166212 180100 166276 180164
rect 335676 180100 335740 180164
rect 160692 179964 160756 180028
rect 346348 179344 346412 179348
rect 346348 179288 346362 179344
rect 346362 179288 346412 179344
rect 346348 179284 346412 179288
rect 342300 179148 342364 179212
rect 249012 178876 249076 178940
rect 259684 178740 259748 178804
rect 256924 178604 256988 178668
rect 332732 178604 332796 178668
rect 110644 178196 110708 178260
rect 167684 178196 167748 178260
rect 166212 178060 166276 178124
rect 97028 177924 97092 177988
rect 99420 177516 99484 177580
rect 101996 177576 102060 177580
rect 101996 177520 102046 177576
rect 102046 177520 102060 177576
rect 101996 177516 102060 177520
rect 104572 177516 104636 177580
rect 106044 177516 106108 177580
rect 113220 177516 113284 177580
rect 118372 177576 118436 177580
rect 118372 177520 118422 177576
rect 118422 177520 118436 177576
rect 118372 177516 118436 177520
rect 121868 177516 121932 177580
rect 124444 177516 124508 177580
rect 131988 177516 132052 177580
rect 133092 177516 133156 177580
rect 249196 177516 249260 177580
rect 318012 177516 318076 177580
rect 334020 177380 334084 177444
rect 52500 177304 52564 177308
rect 52500 177248 52550 177304
rect 52550 177248 52564 177304
rect 52500 177244 52564 177248
rect 336964 177244 337028 177308
rect 114140 176972 114204 177036
rect 120764 176972 120828 177036
rect 122972 177032 123036 177036
rect 122972 176976 123022 177032
rect 123022 176976 123036 177032
rect 122972 176972 123036 176976
rect 103284 176836 103348 176900
rect 167500 176836 167564 176900
rect 106964 176760 107028 176764
rect 106964 176704 107014 176760
rect 107014 176704 107028 176760
rect 106964 176700 107028 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 109540 176700 109604 176764
rect 112116 176700 112180 176764
rect 125732 176760 125796 176764
rect 125732 176704 125782 176760
rect 125782 176704 125796 176760
rect 125732 176700 125796 176704
rect 127020 176760 127084 176764
rect 127020 176704 127070 176760
rect 127070 176704 127084 176760
rect 127020 176700 127084 176704
rect 130700 176760 130764 176764
rect 130700 176704 130750 176760
rect 130750 176704 130764 176760
rect 130700 176700 130764 176704
rect 134380 176760 134444 176764
rect 134380 176704 134430 176760
rect 134430 176704 134444 176760
rect 134380 176700 134444 176704
rect 135668 176760 135732 176764
rect 135668 176704 135718 176760
rect 135718 176704 135732 176760
rect 135668 176700 135732 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 158852 176700 158916 176764
rect 128124 176428 128188 176492
rect 321508 176156 321572 176220
rect 262260 176020 262324 176084
rect 306972 175672 307036 175676
rect 306972 175616 307022 175672
rect 307022 175616 307036 175672
rect 306972 175612 307036 175616
rect 98316 175400 98380 175404
rect 98316 175344 98366 175400
rect 98366 175344 98380 175400
rect 98316 175340 98380 175344
rect 100708 175400 100772 175404
rect 100708 175344 100758 175400
rect 100758 175344 100772 175400
rect 100708 175340 100772 175344
rect 116900 175400 116964 175404
rect 116900 175344 116950 175400
rect 116950 175344 116964 175400
rect 116900 175340 116964 175344
rect 129412 175400 129476 175404
rect 129412 175344 129462 175400
rect 129462 175344 129476 175400
rect 129412 175340 129476 175344
rect 115726 174992 115790 174996
rect 115726 174936 115754 174992
rect 115754 174936 115790 174992
rect 115726 174932 115790 174936
rect 119398 174992 119462 174996
rect 119398 174936 119434 174992
rect 119434 174936 119462 174992
rect 119398 174932 119462 174936
rect 249196 174252 249260 174316
rect 260972 173904 261036 173908
rect 260972 173848 261022 173904
rect 261022 173848 261036 173904
rect 260972 173844 261036 173848
rect 249380 173300 249444 173364
rect 321508 172076 321572 172140
rect 261340 171396 261404 171460
rect 265204 170852 265268 170916
rect 256740 169824 256804 169828
rect 256740 169768 256790 169824
rect 256790 169768 256804 169824
rect 256740 169764 256804 169768
rect 321324 169764 321388 169828
rect 265020 168132 265084 168196
rect 334020 165684 334084 165748
rect 266308 164732 266372 164796
rect 256924 164188 256988 164252
rect 166396 163100 166460 163164
rect 263732 163372 263796 163436
rect 167684 161468 167748 161532
rect 345060 161468 345124 161532
rect 335676 160108 335740 160172
rect 167500 157388 167564 157452
rect 262260 157796 262324 157860
rect 252508 155348 252572 155412
rect 166212 154532 166276 154596
rect 322060 150316 322124 150380
rect 255452 147868 255516 147932
rect 257844 146236 257908 146300
rect 167500 143652 167564 143716
rect 329788 143516 329852 143580
rect 260972 142700 261036 142764
rect 263548 142156 263612 142220
rect 328684 142156 328748 142220
rect 328500 142020 328564 142084
rect 261340 141476 261404 141540
rect 259684 141204 259748 141268
rect 251772 141068 251836 141132
rect 336964 140796 337028 140860
rect 306972 139980 307036 140044
rect 255268 139844 255332 139908
rect 261340 139708 261404 139772
rect 305500 139436 305564 139500
rect 346348 139436 346412 139500
rect 327028 139300 327092 139364
rect 259500 138892 259564 138956
rect 300164 135220 300228 135284
rect 342300 135220 342364 135284
rect 170260 133860 170324 133924
rect 167684 132772 167748 132836
rect 327580 132092 327644 132156
rect 331260 131684 331324 131748
rect 166212 131140 166276 131204
rect 291700 130052 291764 130116
rect 169156 128556 169220 128620
rect 307156 128012 307220 128076
rect 293172 125836 293236 125900
rect 332732 123252 332796 123316
rect 295932 117540 295996 117604
rect 335676 116044 335740 116108
rect 338252 115908 338316 115972
rect 251956 115092 252020 115156
rect 275140 113460 275204 113524
rect 251772 113052 251836 113116
rect 336780 109108 336844 109172
rect 305684 101220 305748 101284
rect 302740 101084 302804 101148
rect 301636 99996 301700 100060
rect 251956 97956 252020 98020
rect 261340 97548 261404 97612
rect 166396 97140 166460 97204
rect 250116 97004 250180 97068
rect 306972 97004 307036 97068
rect 171732 95916 171796 95980
rect 109062 94752 109126 94756
rect 109062 94696 109094 94752
rect 109094 94696 109126 94752
rect 109062 94692 109126 94696
rect 113686 94752 113750 94756
rect 113686 94696 113730 94752
rect 113730 94696 113750 94752
rect 113686 94692 113750 94696
rect 131910 94752 131974 94756
rect 131910 94696 131946 94752
rect 131946 94696 131974 94752
rect 131910 94692 131974 94696
rect 151766 94752 151830 94756
rect 151766 94696 151782 94752
rect 151782 94696 151830 94752
rect 151766 94692 151830 94696
rect 151902 94752 151966 94756
rect 151902 94696 151910 94752
rect 151910 94696 151966 94752
rect 151902 94692 151966 94696
rect 114324 93876 114388 93940
rect 108068 93740 108132 93804
rect 167684 93740 167748 93804
rect 173572 93740 173636 93804
rect 121684 93664 121748 93668
rect 121684 93608 121734 93664
rect 121734 93608 121748 93664
rect 121684 93604 121748 93608
rect 101996 93528 102060 93532
rect 101996 93472 102046 93528
rect 102046 93472 102060 93528
rect 101996 93468 102060 93472
rect 107700 93528 107764 93532
rect 107700 93472 107750 93528
rect 107750 93472 107764 93528
rect 107700 93468 107764 93472
rect 124444 93528 124508 93532
rect 124444 93472 124494 93528
rect 124494 93472 124508 93528
rect 124444 93468 124508 93472
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 119292 93256 119356 93260
rect 119292 93200 119342 93256
rect 119342 93200 119356 93256
rect 119292 93196 119356 93200
rect 74764 92440 74828 92444
rect 74764 92384 74814 92440
rect 74814 92384 74828 92440
rect 74764 92380 74828 92384
rect 85620 92380 85684 92444
rect 93900 92380 93964 92444
rect 101812 92440 101876 92444
rect 101812 92384 101862 92440
rect 101862 92384 101876 92440
rect 101812 92380 101876 92384
rect 115060 92380 115124 92444
rect 115428 92440 115492 92444
rect 115428 92384 115478 92440
rect 115478 92384 115492 92440
rect 115428 92380 115492 92384
rect 120212 92380 120276 92444
rect 124076 92440 124140 92444
rect 124076 92384 124126 92440
rect 124126 92384 124140 92440
rect 124076 92380 124140 92384
rect 125916 92440 125980 92444
rect 125916 92384 125966 92440
rect 125966 92384 125980 92440
rect 125916 92380 125980 92384
rect 133092 92440 133156 92444
rect 133092 92384 133142 92440
rect 133142 92384 133156 92440
rect 133092 92380 133156 92384
rect 151676 92440 151740 92444
rect 151676 92384 151726 92440
rect 151726 92384 151740 92440
rect 151676 92380 151740 92384
rect 174492 92380 174556 92444
rect 111932 92244 111996 92308
rect 166396 92244 166460 92308
rect 106044 92108 106108 92172
rect 88932 91700 88996 91764
rect 112300 91760 112364 91764
rect 112300 91704 112350 91760
rect 112350 91704 112364 91760
rect 112300 91700 112364 91704
rect 122972 91700 123036 91764
rect 151308 91700 151372 91764
rect 104204 91564 104268 91628
rect 106780 91564 106844 91628
rect 126468 91564 126532 91628
rect 98500 91428 98564 91492
rect 122788 91488 122852 91492
rect 122788 91432 122838 91488
rect 122838 91432 122852 91488
rect 122788 91428 122852 91432
rect 97028 91292 97092 91356
rect 98132 91292 98196 91356
rect 118188 91352 118252 91356
rect 118188 91296 118238 91352
rect 118238 91296 118252 91352
rect 118188 91292 118252 91296
rect 84332 91156 84396 91220
rect 86724 91216 86788 91220
rect 86724 91160 86774 91216
rect 86774 91160 86788 91216
rect 86724 91156 86788 91160
rect 87092 91156 87156 91220
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91216 95068 91220
rect 95004 91160 95054 91216
rect 95054 91160 95068 91216
rect 95004 91156 95068 91160
rect 96108 91156 96172 91220
rect 97212 91156 97276 91220
rect 99236 91216 99300 91220
rect 99236 91160 99250 91216
rect 99250 91160 99300 91216
rect 99236 91156 99300 91160
rect 99604 91156 99668 91220
rect 100524 91156 100588 91220
rect 101628 91156 101692 91220
rect 102916 91216 102980 91220
rect 102916 91160 102966 91216
rect 102966 91160 102980 91216
rect 102916 91156 102980 91160
rect 103284 91156 103348 91220
rect 104572 91216 104636 91220
rect 104572 91160 104622 91216
rect 104622 91160 104636 91216
rect 104572 91156 104636 91160
rect 105124 91156 105188 91220
rect 106412 91156 106476 91220
rect 109540 91156 109604 91220
rect 110644 91216 110708 91220
rect 110644 91160 110694 91216
rect 110694 91160 110708 91216
rect 110644 91156 110708 91160
rect 111196 91156 111260 91220
rect 113220 91156 113284 91220
rect 115796 91216 115860 91220
rect 115796 91160 115810 91216
rect 115810 91160 115860 91216
rect 115796 91156 115860 91160
rect 116716 91216 116780 91220
rect 116716 91160 116766 91216
rect 116766 91160 116780 91216
rect 116716 91156 116780 91160
rect 117084 91216 117148 91220
rect 117084 91160 117134 91216
rect 117134 91160 117148 91216
rect 117084 91156 117148 91160
rect 118004 91156 118068 91220
rect 119660 91156 119724 91220
rect 120580 91156 120644 91220
rect 122052 91156 122116 91220
rect 125364 91156 125428 91220
rect 126652 91156 126716 91220
rect 127572 91156 127636 91220
rect 129412 91156 129476 91220
rect 130700 91156 130764 91220
rect 134380 91156 134444 91220
rect 135668 91156 135732 91220
rect 167500 91020 167564 91084
rect 307156 89116 307220 89180
rect 178908 88980 178972 89044
rect 166212 86804 166276 86868
rect 170260 84084 170324 84148
rect 179644 79324 179708 79388
rect 169156 78508 169220 78572
rect 300164 69532 300228 69596
rect 301636 62732 301700 62796
rect 293172 59876 293236 59940
rect 291700 58516 291764 58580
rect 177068 50220 177132 50284
rect 302740 48860 302804 48924
rect 176332 39204 176396 39268
rect 305500 37844 305564 37908
rect 295932 26828 295996 26892
rect 179276 21252 179340 21316
rect 184796 18668 184860 18732
rect 275140 18532 275204 18596
rect 250116 16492 250180 16556
rect 305684 12956 305748 13020
rect 306972 8876 307036 8940
rect 175044 6156 175108 6220
rect 271092 3980 271156 4044
rect 296484 3980 296548 4044
rect 304212 3980 304276 4044
rect 301452 3572 301516 3636
rect 299980 3436 300044 3500
rect 332548 3436 332612 3500
rect 340828 3436 340892 3500
rect 169708 3300 169772 3364
rect 269620 3300 269684 3364
rect 176516 1940 176580 2004
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 50843 583948 50909 583949
rect 50843 583884 50844 583948
rect 50908 583884 50909 583948
rect 50843 583883 50909 583884
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 49555 469844 49621 469845
rect 49555 469780 49556 469844
rect 49620 469780 49621 469844
rect 49555 469779 49621 469780
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 49558 314805 49618 469779
rect 50846 398173 50906 583883
rect 51294 556954 51914 592398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 58939 582588 59005 582589
rect 58939 582524 58940 582588
rect 59004 582524 59005 582588
rect 58939 582523 59005 582524
rect 57835 579188 57901 579189
rect 57835 579124 57836 579188
rect 57900 579124 57901 579188
rect 57835 579123 57901 579124
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 54339 557564 54405 557565
rect 54339 557500 54340 557564
rect 54404 557500 54405 557564
rect 54339 557499 54405 557500
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 53603 464948 53669 464949
rect 53603 464884 53604 464948
rect 53668 464884 53669 464948
rect 53603 464883 53669 464884
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 53419 430676 53485 430677
rect 53419 430612 53420 430676
rect 53484 430612 53485 430676
rect 53419 430611 53485 430612
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 50843 398172 50909 398173
rect 50843 398108 50844 398172
rect 50908 398108 50909 398172
rect 50843 398107 50909 398108
rect 51294 376954 51914 412398
rect 53422 405653 53482 430611
rect 53419 405652 53485 405653
rect 53419 405588 53420 405652
rect 53484 405588 53485 405652
rect 53419 405587 53485 405588
rect 52499 401708 52565 401709
rect 52499 401644 52500 401708
rect 52564 401644 52565 401708
rect 52499 401643 52565 401644
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 49555 314804 49621 314805
rect 49555 314740 49556 314804
rect 49620 314740 49621 314804
rect 49555 314739 49621 314740
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 52502 177309 52562 401643
rect 53606 354653 53666 464883
rect 53603 354652 53669 354653
rect 53603 354588 53604 354652
rect 53668 354588 53669 354652
rect 53603 354587 53669 354588
rect 54342 284341 54402 557499
rect 55627 532268 55693 532269
rect 55627 532204 55628 532268
rect 55692 532204 55693 532268
rect 55627 532203 55693 532204
rect 54339 284340 54405 284341
rect 54339 284276 54340 284340
rect 54404 284276 54405 284340
rect 54339 284275 54405 284276
rect 55630 271829 55690 532203
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 57651 434620 57717 434621
rect 57651 434556 57652 434620
rect 57716 434556 57717 434620
rect 57651 434555 57717 434556
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 57654 404973 57714 434555
rect 57651 404972 57717 404973
rect 57651 404908 57652 404972
rect 57716 404908 57717 404972
rect 57651 404907 57717 404908
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55627 271828 55693 271829
rect 55627 271764 55628 271828
rect 55692 271764 55693 271828
rect 55627 271763 55693 271764
rect 55794 237454 56414 272898
rect 57838 238645 57898 579123
rect 58942 399533 59002 582523
rect 60043 575788 60109 575789
rect 60043 575724 60044 575788
rect 60108 575724 60109 575788
rect 60043 575723 60109 575724
rect 59123 525468 59189 525469
rect 59123 525404 59124 525468
rect 59188 525404 59189 525468
rect 59123 525403 59189 525404
rect 58939 399532 59005 399533
rect 58939 399468 58940 399532
rect 59004 399468 59005 399532
rect 58939 399467 59005 399468
rect 59126 327725 59186 525403
rect 60046 387021 60106 575723
rect 60294 565954 60914 601398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 587000 65414 605898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 587000 69914 610398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 587000 74414 614898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 587000 78914 619398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 587000 83414 587898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 587000 87914 592398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 587000 92414 596898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 587000 96914 601398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 587000 101414 605898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 587000 105914 610398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 587000 110414 614898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 587000 114914 619398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 587000 119414 587898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 587000 123914 592398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 587000 128414 596898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 587000 132914 601398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 587000 137414 605898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 587000 141914 610398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 587000 146414 614898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 587000 150914 619398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 587000 155414 587898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 587000 159914 592398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 587000 164414 596898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 587000 168914 601398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 587000 173414 605898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 587000 177914 610398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 587000 182414 614898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 587000 186914 619398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 587000 191414 587898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 587000 195914 592398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 587000 200414 596898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 587000 204914 601398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 587000 209414 605898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 587000 213914 610398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 587000 218414 614898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 587000 222914 619398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 587000 227414 587898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 587000 231914 592398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 587000 236414 596898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 587000 240914 601398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 587000 245414 605898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 243491 586532 243557 586533
rect 243491 586468 243492 586532
rect 243556 586468 243557 586532
rect 243491 586467 243557 586468
rect 63539 584628 63605 584629
rect 63539 584564 63540 584628
rect 63604 584564 63605 584628
rect 63539 584563 63605 584564
rect 61883 572388 61949 572389
rect 61883 572324 61884 572388
rect 61948 572324 61949 572388
rect 61883 572323 61949 572324
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60043 387020 60109 387021
rect 60043 386956 60044 387020
rect 60108 386956 60109 387020
rect 60043 386955 60109 386956
rect 60294 385954 60914 421398
rect 61886 404429 61946 572323
rect 63542 558245 63602 584563
rect 243307 579596 243373 579597
rect 243307 579532 243308 579596
rect 243372 579532 243373 579596
rect 243307 579531 243373 579532
rect 68208 579454 68528 579486
rect 68208 579218 68250 579454
rect 68486 579218 68528 579454
rect 68208 579134 68528 579218
rect 68208 578898 68250 579134
rect 68486 578898 68528 579134
rect 68208 578866 68528 578898
rect 98928 579454 99248 579486
rect 98928 579218 98970 579454
rect 99206 579218 99248 579454
rect 98928 579134 99248 579218
rect 98928 578898 98970 579134
rect 99206 578898 99248 579134
rect 98928 578866 99248 578898
rect 129648 579454 129968 579486
rect 129648 579218 129690 579454
rect 129926 579218 129968 579454
rect 129648 579134 129968 579218
rect 129648 578898 129690 579134
rect 129926 578898 129968 579134
rect 129648 578866 129968 578898
rect 160368 579454 160688 579486
rect 160368 579218 160410 579454
rect 160646 579218 160688 579454
rect 160368 579134 160688 579218
rect 160368 578898 160410 579134
rect 160646 578898 160688 579134
rect 160368 578866 160688 578898
rect 191088 579454 191408 579486
rect 191088 579218 191130 579454
rect 191366 579218 191408 579454
rect 191088 579134 191408 579218
rect 191088 578898 191130 579134
rect 191366 578898 191408 579134
rect 191088 578866 191408 578898
rect 221808 579454 222128 579486
rect 221808 579218 221850 579454
rect 222086 579218 222128 579454
rect 221808 579134 222128 579218
rect 221808 578898 221850 579134
rect 222086 578898 222128 579134
rect 221808 578866 222128 578898
rect 243310 567210 243370 579531
rect 243494 578917 243554 586467
rect 247171 585444 247237 585445
rect 247171 585380 247172 585444
rect 247236 585380 247237 585444
rect 247171 585379 247237 585380
rect 243675 585172 243741 585173
rect 243675 585108 243676 585172
rect 243740 585108 243741 585172
rect 243675 585107 243741 585108
rect 243678 580957 243738 585107
rect 243675 580956 243741 580957
rect 243675 580892 243676 580956
rect 243740 580892 243741 580956
rect 243675 580891 243741 580892
rect 243491 578916 243557 578917
rect 243491 578852 243492 578916
rect 243556 578852 243557 578916
rect 243491 578851 243557 578852
rect 246987 569668 247053 569669
rect 246987 569604 246988 569668
rect 247052 569604 247053 569668
rect 246987 569603 247053 569604
rect 242942 567150 243370 567210
rect 63539 558244 63605 558245
rect 63539 558180 63540 558244
rect 63604 558180 63605 558244
rect 63539 558179 63605 558180
rect 83568 547954 83888 547986
rect 83568 547718 83610 547954
rect 83846 547718 83888 547954
rect 83568 547634 83888 547718
rect 83568 547398 83610 547634
rect 83846 547398 83888 547634
rect 83568 547366 83888 547398
rect 114288 547954 114608 547986
rect 114288 547718 114330 547954
rect 114566 547718 114608 547954
rect 114288 547634 114608 547718
rect 114288 547398 114330 547634
rect 114566 547398 114608 547634
rect 114288 547366 114608 547398
rect 145008 547954 145328 547986
rect 145008 547718 145050 547954
rect 145286 547718 145328 547954
rect 145008 547634 145328 547718
rect 145008 547398 145050 547634
rect 145286 547398 145328 547634
rect 145008 547366 145328 547398
rect 175728 547954 176048 547986
rect 175728 547718 175770 547954
rect 176006 547718 176048 547954
rect 175728 547634 176048 547718
rect 175728 547398 175770 547634
rect 176006 547398 176048 547634
rect 175728 547366 176048 547398
rect 206448 547954 206768 547986
rect 206448 547718 206490 547954
rect 206726 547718 206768 547954
rect 206448 547634 206768 547718
rect 206448 547398 206490 547634
rect 206726 547398 206768 547634
rect 206448 547366 206768 547398
rect 237168 547954 237488 547986
rect 237168 547718 237210 547954
rect 237446 547718 237488 547954
rect 237168 547634 237488 547718
rect 237168 547398 237210 547634
rect 237446 547398 237488 547634
rect 237168 547366 237488 547398
rect 68208 543454 68528 543486
rect 68208 543218 68250 543454
rect 68486 543218 68528 543454
rect 68208 543134 68528 543218
rect 68208 542898 68250 543134
rect 68486 542898 68528 543134
rect 68208 542866 68528 542898
rect 98928 543454 99248 543486
rect 98928 543218 98970 543454
rect 99206 543218 99248 543454
rect 98928 543134 99248 543218
rect 98928 542898 98970 543134
rect 99206 542898 99248 543134
rect 98928 542866 99248 542898
rect 129648 543454 129968 543486
rect 129648 543218 129690 543454
rect 129926 543218 129968 543454
rect 129648 543134 129968 543218
rect 129648 542898 129690 543134
rect 129926 542898 129968 543134
rect 129648 542866 129968 542898
rect 160368 543454 160688 543486
rect 160368 543218 160410 543454
rect 160646 543218 160688 543454
rect 160368 543134 160688 543218
rect 160368 542898 160410 543134
rect 160646 542898 160688 543134
rect 160368 542866 160688 542898
rect 191088 543454 191408 543486
rect 191088 543218 191130 543454
rect 191366 543218 191408 543454
rect 191088 543134 191408 543218
rect 191088 542898 191130 543134
rect 191366 542898 191408 543134
rect 191088 542866 191408 542898
rect 221808 543454 222128 543486
rect 221808 543218 221850 543454
rect 222086 543218 222128 543454
rect 221808 543134 222128 543218
rect 221808 542898 221850 543134
rect 222086 542898 222128 543134
rect 221808 542866 222128 542898
rect 83568 511954 83888 511986
rect 63539 511868 63605 511869
rect 63539 511804 63540 511868
rect 63604 511804 63605 511868
rect 63539 511803 63605 511804
rect 62067 510508 62133 510509
rect 62067 510444 62068 510508
rect 62132 510444 62133 510508
rect 62067 510443 62133 510444
rect 62070 485893 62130 510443
rect 62067 485892 62133 485893
rect 62067 485828 62068 485892
rect 62132 485828 62133 485892
rect 62067 485827 62133 485828
rect 63355 448628 63421 448629
rect 63355 448564 63356 448628
rect 63420 448564 63421 448628
rect 63355 448563 63421 448564
rect 63171 421428 63237 421429
rect 63171 421364 63172 421428
rect 63236 421364 63237 421428
rect 63171 421363 63237 421364
rect 63174 404565 63234 421363
rect 63171 404564 63237 404565
rect 63171 404500 63172 404564
rect 63236 404500 63237 404564
rect 63171 404499 63237 404500
rect 61883 404428 61949 404429
rect 61883 404364 61884 404428
rect 61948 404364 61949 404428
rect 61883 404363 61949 404364
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 59123 327724 59189 327725
rect 59123 327660 59124 327724
rect 59188 327660 59189 327724
rect 59123 327659 59189 327660
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 63171 254012 63237 254013
rect 63171 253948 63172 254012
rect 63236 253948 63237 254012
rect 63171 253947 63237 253948
rect 61883 244492 61949 244493
rect 61883 244428 61884 244492
rect 61948 244428 61949 244492
rect 61883 244427 61949 244428
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 57835 238644 57901 238645
rect 57835 238580 57836 238644
rect 57900 238580 57901 238644
rect 57835 238579 57901 238580
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 52499 177308 52565 177309
rect 52499 177244 52500 177308
rect 52564 177244 52565 177308
rect 52499 177243 52565 177244
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 241398
rect 61886 237285 61946 244427
rect 61883 237284 61949 237285
rect 61883 237220 61884 237284
rect 61948 237220 61949 237284
rect 61883 237219 61949 237220
rect 63174 222189 63234 253947
rect 63358 252517 63418 448563
rect 63542 398037 63602 511803
rect 83568 511718 83610 511954
rect 83846 511718 83888 511954
rect 83568 511634 83888 511718
rect 83568 511398 83610 511634
rect 83846 511398 83888 511634
rect 83568 511366 83888 511398
rect 114288 511954 114608 511986
rect 114288 511718 114330 511954
rect 114566 511718 114608 511954
rect 114288 511634 114608 511718
rect 114288 511398 114330 511634
rect 114566 511398 114608 511634
rect 114288 511366 114608 511398
rect 145008 511954 145328 511986
rect 145008 511718 145050 511954
rect 145286 511718 145328 511954
rect 145008 511634 145328 511718
rect 145008 511398 145050 511634
rect 145286 511398 145328 511634
rect 145008 511366 145328 511398
rect 175728 511954 176048 511986
rect 175728 511718 175770 511954
rect 176006 511718 176048 511954
rect 175728 511634 176048 511718
rect 175728 511398 175770 511634
rect 176006 511398 176048 511634
rect 175728 511366 176048 511398
rect 206448 511954 206768 511986
rect 206448 511718 206490 511954
rect 206726 511718 206768 511954
rect 206448 511634 206768 511718
rect 206448 511398 206490 511634
rect 206726 511398 206768 511634
rect 206448 511366 206768 511398
rect 237168 511954 237488 511986
rect 237168 511718 237210 511954
rect 237446 511718 237488 511954
rect 237168 511634 237488 511718
rect 237168 511398 237210 511634
rect 237446 511398 237488 511634
rect 237168 511366 237488 511398
rect 68208 507454 68528 507486
rect 68208 507218 68250 507454
rect 68486 507218 68528 507454
rect 68208 507134 68528 507218
rect 68208 506898 68250 507134
rect 68486 506898 68528 507134
rect 68208 506866 68528 506898
rect 98928 507454 99248 507486
rect 98928 507218 98970 507454
rect 99206 507218 99248 507454
rect 98928 507134 99248 507218
rect 98928 506898 98970 507134
rect 99206 506898 99248 507134
rect 98928 506866 99248 506898
rect 129648 507454 129968 507486
rect 129648 507218 129690 507454
rect 129926 507218 129968 507454
rect 129648 507134 129968 507218
rect 129648 506898 129690 507134
rect 129926 506898 129968 507134
rect 129648 506866 129968 506898
rect 160368 507454 160688 507486
rect 160368 507218 160410 507454
rect 160646 507218 160688 507454
rect 160368 507134 160688 507218
rect 160368 506898 160410 507134
rect 160646 506898 160688 507134
rect 160368 506866 160688 506898
rect 191088 507454 191408 507486
rect 191088 507218 191130 507454
rect 191366 507218 191408 507454
rect 191088 507134 191408 507218
rect 191088 506898 191130 507134
rect 191366 506898 191408 507134
rect 191088 506866 191408 506898
rect 221808 507454 222128 507486
rect 221808 507218 221850 507454
rect 222086 507218 222128 507454
rect 221808 507134 222128 507218
rect 221808 506898 221850 507134
rect 222086 506898 222128 507134
rect 221808 506866 222128 506898
rect 83568 475954 83888 475986
rect 83568 475718 83610 475954
rect 83846 475718 83888 475954
rect 83568 475634 83888 475718
rect 83568 475398 83610 475634
rect 83846 475398 83888 475634
rect 83568 475366 83888 475398
rect 114288 475954 114608 475986
rect 114288 475718 114330 475954
rect 114566 475718 114608 475954
rect 114288 475634 114608 475718
rect 114288 475398 114330 475634
rect 114566 475398 114608 475634
rect 114288 475366 114608 475398
rect 145008 475954 145328 475986
rect 145008 475718 145050 475954
rect 145286 475718 145328 475954
rect 145008 475634 145328 475718
rect 145008 475398 145050 475634
rect 145286 475398 145328 475634
rect 145008 475366 145328 475398
rect 175728 475954 176048 475986
rect 175728 475718 175770 475954
rect 176006 475718 176048 475954
rect 175728 475634 176048 475718
rect 175728 475398 175770 475634
rect 176006 475398 176048 475634
rect 175728 475366 176048 475398
rect 206448 475954 206768 475986
rect 206448 475718 206490 475954
rect 206726 475718 206768 475954
rect 206448 475634 206768 475718
rect 206448 475398 206490 475634
rect 206726 475398 206768 475634
rect 206448 475366 206768 475398
rect 237168 475954 237488 475986
rect 237168 475718 237210 475954
rect 237446 475718 237488 475954
rect 237168 475634 237488 475718
rect 237168 475398 237210 475634
rect 237446 475398 237488 475634
rect 237168 475366 237488 475398
rect 63723 473244 63789 473245
rect 63723 473180 63724 473244
rect 63788 473180 63789 473244
rect 63723 473179 63789 473180
rect 63726 449989 63786 473179
rect 68208 471454 68528 471486
rect 68208 471218 68250 471454
rect 68486 471218 68528 471454
rect 68208 471134 68528 471218
rect 68208 470898 68250 471134
rect 68486 470898 68528 471134
rect 68208 470866 68528 470898
rect 98928 471454 99248 471486
rect 98928 471218 98970 471454
rect 99206 471218 99248 471454
rect 98928 471134 99248 471218
rect 98928 470898 98970 471134
rect 99206 470898 99248 471134
rect 98928 470866 99248 470898
rect 129648 471454 129968 471486
rect 129648 471218 129690 471454
rect 129926 471218 129968 471454
rect 129648 471134 129968 471218
rect 129648 470898 129690 471134
rect 129926 470898 129968 471134
rect 129648 470866 129968 470898
rect 160368 471454 160688 471486
rect 160368 471218 160410 471454
rect 160646 471218 160688 471454
rect 160368 471134 160688 471218
rect 160368 470898 160410 471134
rect 160646 470898 160688 471134
rect 160368 470866 160688 470898
rect 191088 471454 191408 471486
rect 191088 471218 191130 471454
rect 191366 471218 191408 471454
rect 191088 471134 191408 471218
rect 191088 470898 191130 471134
rect 191366 470898 191408 471134
rect 191088 470866 191408 470898
rect 221808 471454 222128 471486
rect 221808 471218 221850 471454
rect 222086 471218 222128 471454
rect 221808 471134 222128 471218
rect 221808 470898 221850 471134
rect 222086 470898 222128 471134
rect 221808 470866 222128 470898
rect 63723 449988 63789 449989
rect 63723 449924 63724 449988
rect 63788 449924 63789 449988
rect 63723 449923 63789 449924
rect 83568 439954 83888 439986
rect 83568 439718 83610 439954
rect 83846 439718 83888 439954
rect 83568 439634 83888 439718
rect 83568 439398 83610 439634
rect 83846 439398 83888 439634
rect 83568 439366 83888 439398
rect 114288 439954 114608 439986
rect 114288 439718 114330 439954
rect 114566 439718 114608 439954
rect 114288 439634 114608 439718
rect 114288 439398 114330 439634
rect 114566 439398 114608 439634
rect 114288 439366 114608 439398
rect 145008 439954 145328 439986
rect 145008 439718 145050 439954
rect 145286 439718 145328 439954
rect 145008 439634 145328 439718
rect 145008 439398 145050 439634
rect 145286 439398 145328 439634
rect 145008 439366 145328 439398
rect 175728 439954 176048 439986
rect 175728 439718 175770 439954
rect 176006 439718 176048 439954
rect 175728 439634 176048 439718
rect 175728 439398 175770 439634
rect 176006 439398 176048 439634
rect 175728 439366 176048 439398
rect 206448 439954 206768 439986
rect 206448 439718 206490 439954
rect 206726 439718 206768 439954
rect 206448 439634 206768 439718
rect 206448 439398 206490 439634
rect 206726 439398 206768 439634
rect 206448 439366 206768 439398
rect 237168 439954 237488 439986
rect 237168 439718 237210 439954
rect 237446 439718 237488 439954
rect 237168 439634 237488 439718
rect 237168 439398 237210 439634
rect 237446 439398 237488 439634
rect 237168 439366 237488 439398
rect 68208 435454 68528 435486
rect 68208 435218 68250 435454
rect 68486 435218 68528 435454
rect 68208 435134 68528 435218
rect 68208 434898 68250 435134
rect 68486 434898 68528 435134
rect 68208 434866 68528 434898
rect 98928 435454 99248 435486
rect 98928 435218 98970 435454
rect 99206 435218 99248 435454
rect 98928 435134 99248 435218
rect 98928 434898 98970 435134
rect 99206 434898 99248 435134
rect 98928 434866 99248 434898
rect 129648 435454 129968 435486
rect 129648 435218 129690 435454
rect 129926 435218 129968 435454
rect 129648 435134 129968 435218
rect 129648 434898 129690 435134
rect 129926 434898 129968 435134
rect 129648 434866 129968 434898
rect 160368 435454 160688 435486
rect 160368 435218 160410 435454
rect 160646 435218 160688 435454
rect 160368 435134 160688 435218
rect 160368 434898 160410 435134
rect 160646 434898 160688 435134
rect 160368 434866 160688 434898
rect 191088 435454 191408 435486
rect 191088 435218 191130 435454
rect 191366 435218 191408 435454
rect 191088 435134 191408 435218
rect 191088 434898 191130 435134
rect 191366 434898 191408 435134
rect 191088 434866 191408 434898
rect 221808 435454 222128 435486
rect 221808 435218 221850 435454
rect 222086 435218 222128 435454
rect 221808 435134 222128 435218
rect 221808 434898 221850 435134
rect 222086 434898 222128 435134
rect 221808 434866 222128 434898
rect 64091 429316 64157 429317
rect 64091 429252 64092 429316
rect 64156 429252 64157 429316
rect 64091 429251 64157 429252
rect 63539 398036 63605 398037
rect 63539 397972 63540 398036
rect 63604 397972 63605 398036
rect 63539 397971 63605 397972
rect 64094 356693 64154 429251
rect 66851 403748 66917 403749
rect 66851 403684 66852 403748
rect 66916 403684 66917 403748
rect 66851 403683 66917 403684
rect 64794 390454 65414 403000
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64091 356692 64157 356693
rect 64091 356628 64092 356692
rect 64156 356628 64157 356692
rect 64091 356627 64157 356628
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64643 294540 64709 294541
rect 64643 294476 64644 294540
rect 64708 294476 64709 294540
rect 64643 294475 64709 294476
rect 64459 256868 64525 256869
rect 64459 256804 64460 256868
rect 64524 256804 64525 256868
rect 64459 256803 64525 256804
rect 63355 252516 63421 252517
rect 63355 252452 63356 252516
rect 63420 252452 63421 252516
rect 63355 252451 63421 252452
rect 64462 235245 64522 256803
rect 64459 235244 64525 235245
rect 64459 235180 64460 235244
rect 64524 235180 64525 235244
rect 64459 235179 64525 235180
rect 63171 222188 63237 222189
rect 63171 222124 63172 222188
rect 63236 222124 63237 222188
rect 63171 222123 63237 222124
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 64646 200701 64706 294475
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 66854 253061 66914 403683
rect 69294 394954 69914 403000
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 73794 399454 74414 403000
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 70899 378180 70965 378181
rect 70899 378116 70900 378180
rect 70964 378116 70965 378180
rect 70899 378115 70965 378116
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69059 298756 69125 298757
rect 69059 298692 69060 298756
rect 69124 298692 69125 298756
rect 69059 298691 69125 298692
rect 66851 253060 66917 253061
rect 66851 252996 66852 253060
rect 66916 252996 66917 253060
rect 66851 252995 66917 252996
rect 67403 253060 67469 253061
rect 67403 252996 67404 253060
rect 67468 252996 67469 253060
rect 67403 252995 67469 252996
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64643 200700 64709 200701
rect 64643 200636 64644 200700
rect 64708 200636 64709 200700
rect 64643 200635 64709 200636
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 174454 65414 209898
rect 67406 193901 67466 252995
rect 69062 252381 69122 298691
rect 69294 294000 69914 322398
rect 70902 296730 70962 378115
rect 70534 296670 70962 296730
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 70534 288149 70594 296670
rect 73794 294000 74414 326898
rect 78294 367954 78914 403000
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 294000 78914 295398
rect 82794 372454 83414 403000
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 294000 83414 299898
rect 87294 376954 87914 403000
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 294000 87914 304398
rect 91794 381454 92414 403000
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 96294 385954 96914 403000
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 294000 96914 313398
rect 100794 390454 101414 403000
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 294000 101414 317898
rect 105294 394954 105914 403000
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 294000 105914 322398
rect 109794 399454 110414 403000
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 114294 367954 114914 403000
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 294000 114914 295398
rect 118794 372454 119414 403000
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 123294 376954 123914 403000
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 119659 359412 119725 359413
rect 119659 359348 119660 359412
rect 119724 359348 119725 359412
rect 119659 359347 119725 359348
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 294000 119414 299898
rect 70531 288148 70597 288149
rect 70531 288084 70532 288148
rect 70596 288084 70597 288148
rect 70531 288083 70597 288084
rect 119662 283389 119722 359347
rect 123294 340954 123914 376398
rect 127794 381454 128414 403000
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 132294 385954 132914 403000
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 129043 357644 129109 357645
rect 129043 357580 129044 357644
rect 129108 357580 129109 357644
rect 129043 357579 129109 357580
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 125731 341460 125797 341461
rect 125731 341396 125732 341460
rect 125796 341396 125797 341460
rect 125731 341395 125797 341396
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 122051 292636 122117 292637
rect 122051 292572 122052 292636
rect 122116 292572 122117 292636
rect 122051 292571 122117 292572
rect 120027 291956 120093 291957
rect 120027 291892 120028 291956
rect 120092 291892 120093 291956
rect 120027 291891 120093 291892
rect 119659 283388 119725 283389
rect 119659 283324 119660 283388
rect 119724 283324 119725 283388
rect 119659 283323 119725 283324
rect 120030 277410 120090 291891
rect 120579 285972 120645 285973
rect 120579 285908 120580 285972
rect 120644 285908 120645 285972
rect 120579 285907 120645 285908
rect 119846 277350 120090 277410
rect 89568 259954 89888 259986
rect 89568 259718 89610 259954
rect 89846 259718 89888 259954
rect 89568 259634 89888 259718
rect 89568 259398 89610 259634
rect 89846 259398 89888 259634
rect 89568 259366 89888 259398
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 69059 252380 69125 252381
rect 69059 252316 69060 252380
rect 69124 252316 69125 252380
rect 69059 252315 69125 252316
rect 69294 214954 69914 238000
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 67403 193900 67469 193901
rect 67403 193836 67404 193900
rect 67468 193836 67469 193900
rect 67403 193835 67469 193836
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 176600 69914 178398
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 78294 223954 78914 238000
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 176600 78914 187398
rect 82794 228454 83414 238000
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 176600 83414 191898
rect 87294 232954 87914 238000
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 176600 87914 196398
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 105294 214954 105914 238000
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 97027 177988 97093 177989
rect 97027 177924 97028 177988
rect 97092 177924 97093 177988
rect 97027 177923 97093 177924
rect 97030 175130 97090 177923
rect 99419 177580 99485 177581
rect 99419 177516 99420 177580
rect 99484 177516 99485 177580
rect 99419 177515 99485 177516
rect 101995 177580 102061 177581
rect 101995 177516 101996 177580
rect 102060 177516 102061 177580
rect 101995 177515 102061 177516
rect 104571 177580 104637 177581
rect 104571 177516 104572 177580
rect 104636 177516 104637 177580
rect 104571 177515 104637 177516
rect 98315 175404 98381 175405
rect 98315 175340 98316 175404
rect 98380 175340 98381 175404
rect 98315 175339 98381 175340
rect 96960 175070 97090 175130
rect 98318 175130 98378 175339
rect 99422 175130 99482 177515
rect 100707 175404 100773 175405
rect 100707 175340 100708 175404
rect 100772 175340 100773 175404
rect 100707 175339 100773 175340
rect 98318 175070 98380 175130
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 175339
rect 101998 175130 102058 177515
rect 103283 176900 103349 176901
rect 103283 176836 103284 176900
rect 103348 176836 103349 176900
rect 103283 176835 103349 176836
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176835
rect 104574 175130 104634 177515
rect 105294 176600 105914 178398
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 106043 177580 106109 177581
rect 106043 177516 106044 177580
rect 106108 177516 106109 177580
rect 106043 177515 106109 177516
rect 106046 175130 106106 177515
rect 106963 176764 107029 176765
rect 106963 176700 106964 176764
rect 107028 176700 107029 176764
rect 106963 176699 107029 176700
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 106106 175130
rect 106966 175130 107026 176699
rect 108070 175130 108130 176699
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 114294 223954 114914 238000
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 110643 178260 110709 178261
rect 110643 178196 110644 178260
rect 110708 178196 110709 178260
rect 110643 178195 110709 178196
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 178195
rect 113219 177580 113285 177581
rect 113219 177516 113220 177580
rect 113284 177516 113285 177580
rect 113219 177515 113285 177516
rect 112115 176764 112181 176765
rect 112115 176700 112116 176764
rect 112180 176700 112181 176764
rect 112115 176699 112181 176700
rect 112118 175130 112178 176699
rect 113222 175130 113282 177515
rect 114139 177036 114205 177037
rect 114139 176972 114140 177036
rect 114204 176972 114205 177036
rect 114139 176971 114205 176972
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114142 175130 114202 176971
rect 114294 176600 114914 187398
rect 118794 228454 119414 238000
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 119846 210357 119906 277350
rect 120582 237149 120642 285907
rect 122054 255917 122114 292571
rect 123294 268954 123914 304398
rect 124259 301476 124325 301477
rect 124259 301412 124260 301476
rect 124324 301412 124325 301476
rect 124259 301411 124325 301412
rect 124075 290460 124141 290461
rect 124075 290396 124076 290460
rect 124140 290396 124141 290460
rect 124075 290395 124141 290396
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 122051 255916 122117 255917
rect 122051 255852 122052 255916
rect 122116 255852 122117 255916
rect 122051 255851 122117 255852
rect 120579 237148 120645 237149
rect 120579 237084 120580 237148
rect 120644 237084 120645 237148
rect 120579 237083 120645 237084
rect 123294 232954 123914 268398
rect 124078 238781 124138 290395
rect 124262 287061 124322 301411
rect 124259 287060 124325 287061
rect 124259 286996 124260 287060
rect 124324 286996 124325 287060
rect 124259 286995 124325 286996
rect 124262 286653 124322 286995
rect 124259 286652 124325 286653
rect 124259 286588 124260 286652
rect 124324 286588 124325 286652
rect 124259 286587 124325 286588
rect 125734 285701 125794 341395
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 125731 285700 125797 285701
rect 125731 285636 125732 285700
rect 125796 285636 125797 285700
rect 125731 285635 125797 285636
rect 126099 283252 126165 283253
rect 126099 283188 126100 283252
rect 126164 283188 126165 283252
rect 126099 283187 126165 283188
rect 126102 241501 126162 283187
rect 127794 273454 128414 308898
rect 128859 305012 128925 305013
rect 128859 304948 128860 305012
rect 128924 304948 128925 305012
rect 128859 304947 128925 304948
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 126099 241500 126165 241501
rect 126099 241436 126100 241500
rect 126164 241436 126165 241500
rect 126099 241435 126165 241436
rect 124075 238780 124141 238781
rect 124075 238716 124076 238780
rect 124140 238716 124141 238780
rect 124075 238715 124141 238716
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 119843 210356 119909 210357
rect 119843 210292 119844 210356
rect 119908 210292 119909 210356
rect 119843 210291 119909 210292
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118371 177580 118437 177581
rect 118371 177516 118372 177580
rect 118436 177516 118437 177580
rect 118371 177515 118437 177516
rect 116899 175404 116965 175405
rect 116899 175340 116900 175404
rect 116964 175340 116965 175404
rect 116899 175339 116965 175340
rect 116902 175130 116962 175339
rect 118374 175130 118434 177515
rect 118794 176600 119414 191898
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 121867 177580 121933 177581
rect 121867 177516 121868 177580
rect 121932 177516 121933 177580
rect 121867 177515 121933 177516
rect 120763 177036 120829 177037
rect 120763 176972 120764 177036
rect 120828 176972 120829 177036
rect 120763 176971 120829 176972
rect 120766 175130 120826 176971
rect 121870 175130 121930 177515
rect 122971 177036 123037 177037
rect 122971 176972 122972 177036
rect 123036 176972 123037 177036
rect 122971 176971 123037 176972
rect 114142 175070 114428 175130
rect 116902 175070 117012 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115725 174996 115791 174997
rect 115725 174932 115726 174996
rect 115790 174932 115791 174996
rect 115725 174931 115791 174932
rect 115728 174494 115788 174931
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 122974 175130 123034 176971
rect 123294 176600 123914 196398
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 128862 202197 128922 304947
rect 129046 289237 129106 357579
rect 132294 349954 132914 385398
rect 136794 390454 137414 403000
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 134379 367164 134445 367165
rect 134379 367100 134380 367164
rect 134444 367100 134445 367164
rect 134379 367099 134445 367100
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 130331 299572 130397 299573
rect 130331 299508 130332 299572
rect 130396 299508 130397 299572
rect 130331 299507 130397 299508
rect 129043 289236 129109 289237
rect 129043 289172 129044 289236
rect 129108 289172 129109 289236
rect 129043 289171 129109 289172
rect 130334 213213 130394 299507
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 130331 213212 130397 213213
rect 130331 213148 130332 213212
rect 130396 213148 130397 213212
rect 130331 213147 130397 213148
rect 132294 205954 132914 241398
rect 134382 237013 134442 367099
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 141294 394954 141914 403000
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 138611 301068 138677 301069
rect 138611 301004 138612 301068
rect 138676 301004 138677 301068
rect 138611 301003 138677 301004
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 134379 237012 134445 237013
rect 134379 236948 134380 237012
rect 134444 236948 134445 237012
rect 134379 236947 134445 236948
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 128859 202196 128925 202197
rect 128859 202132 128860 202196
rect 128924 202132 128925 202196
rect 128859 202131 128925 202132
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 124443 177580 124509 177581
rect 124443 177516 124444 177580
rect 124508 177516 124509 177580
rect 124443 177515 124509 177516
rect 124446 175130 124506 177515
rect 125731 176764 125797 176765
rect 125731 176700 125732 176764
rect 125796 176700 125797 176764
rect 125731 176699 125797 176700
rect 127019 176764 127085 176765
rect 127019 176700 127020 176764
rect 127084 176700 127085 176764
rect 127019 176699 127085 176700
rect 125734 175130 125794 176699
rect 127022 175130 127082 176699
rect 127794 176600 128414 200898
rect 131987 177580 132053 177581
rect 131987 177516 131988 177580
rect 132052 177516 132053 177580
rect 131987 177515 132053 177516
rect 130699 176764 130765 176765
rect 130699 176700 130700 176764
rect 130764 176700 130765 176764
rect 130699 176699 130765 176700
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 129411 175404 129477 175405
rect 129411 175340 129412 175404
rect 129476 175340 129477 175404
rect 129411 175339 129477 175340
rect 122974 175070 123132 175130
rect 118312 174494 118372 175070
rect 119397 174996 119463 174997
rect 119397 174932 119398 174996
rect 119462 174932 119463 174996
rect 119397 174931 119463 174932
rect 119400 174494 119460 174931
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 175339
rect 130702 175130 130762 176699
rect 129414 175070 129524 175130
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 131990 175130 132050 177515
rect 132294 176600 132914 205398
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 133091 177580 133157 177581
rect 133091 177516 133092 177580
rect 133156 177516 133157 177580
rect 133091 177515 133157 177516
rect 133094 175130 133154 177515
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 135667 176764 135733 176765
rect 135667 176700 135668 176764
rect 135732 176700 135733 176764
rect 135667 176699 135733 176700
rect 134382 175130 134442 176699
rect 131990 175070 132108 175130
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135670 175130 135730 176699
rect 136794 176600 137414 209898
rect 138614 196621 138674 301003
rect 141294 286954 141914 322398
rect 145794 399454 146414 403000
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 146891 368524 146957 368525
rect 146891 368460 146892 368524
rect 146956 368460 146957 368524
rect 146891 368459 146957 368460
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 144683 301476 144749 301477
rect 144683 301412 144684 301476
rect 144748 301412 144749 301476
rect 144683 301411 144749 301412
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 144686 243541 144746 301411
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 144683 243540 144749 243541
rect 144683 243476 144684 243540
rect 144748 243476 144749 243540
rect 144683 243475 144749 243476
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 138611 196620 138677 196621
rect 138611 196556 138612 196620
rect 138676 196556 138677 196620
rect 138611 196555 138677 196556
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 176600 141914 178398
rect 145794 219454 146414 254898
rect 146894 242997 146954 368459
rect 150294 367954 150914 403000
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 154794 372454 155414 403000
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 152411 352612 152477 352613
rect 152411 352548 152412 352612
rect 152476 352548 152477 352612
rect 152411 352547 152477 352548
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 148179 303652 148245 303653
rect 148179 303588 148180 303652
rect 148244 303588 148245 303652
rect 148179 303587 148245 303588
rect 146891 242996 146957 242997
rect 146891 242932 146892 242996
rect 146956 242932 146957 242996
rect 146891 242931 146957 242932
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 148182 188325 148242 303587
rect 150294 295954 150914 331398
rect 152414 301205 152474 352547
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 152411 301204 152477 301205
rect 152411 301140 152412 301204
rect 152476 301140 152477 301204
rect 152411 301139 152477 301140
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 149651 272644 149717 272645
rect 149651 272580 149652 272644
rect 149716 272580 149717 272644
rect 149651 272579 149717 272580
rect 149654 265029 149714 272579
rect 149651 265028 149717 265029
rect 149651 264964 149652 265028
rect 149716 264964 149717 265028
rect 149651 264963 149717 264964
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 149651 255916 149717 255917
rect 149651 255852 149652 255916
rect 149716 255852 149717 255916
rect 149651 255851 149717 255852
rect 149654 222053 149714 255851
rect 150294 223954 150914 259398
rect 152414 241773 152474 301139
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 153699 296988 153765 296989
rect 153699 296924 153700 296988
rect 153764 296924 153765 296988
rect 153699 296923 153765 296924
rect 152411 241772 152477 241773
rect 152411 241708 152412 241772
rect 152476 241708 152477 241772
rect 152411 241707 152477 241708
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 149651 222052 149717 222053
rect 149651 221988 149652 222052
rect 149716 221988 149717 222052
rect 149651 221987 149717 221988
rect 148179 188324 148245 188325
rect 148179 188260 148180 188324
rect 148244 188260 148245 188324
rect 148179 188259 148245 188260
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 148182 175130 148242 176699
rect 150294 176600 150914 187398
rect 153702 184245 153762 296923
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 153699 184244 153765 184245
rect 153699 184180 153700 184244
rect 153764 184180 153765 184244
rect 153699 184179 153765 184180
rect 154794 176600 155414 191898
rect 159294 376954 159914 403000
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 163794 381454 164414 403000
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 161979 314804 162045 314805
rect 161979 314740 161980 314804
rect 162044 314740 162045 314804
rect 161979 314739 162045 314740
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 160691 295492 160757 295493
rect 160691 295428 160692 295492
rect 160756 295428 160757 295492
rect 160691 295427 160757 295428
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 159294 176600 159914 196398
rect 160694 180029 160754 295427
rect 161982 238645 162042 314739
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 168294 385954 168914 403000
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 172794 390454 173414 403000
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172283 359412 172349 359413
rect 172283 359348 172284 359412
rect 172348 359348 172349 359412
rect 172283 359347 172349 359348
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 169707 295628 169773 295629
rect 169707 295564 169708 295628
rect 169772 295564 169773 295628
rect 169707 295563 169773 295564
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 166395 276044 166461 276045
rect 166395 275980 166396 276044
rect 166460 275980 166461 276044
rect 166395 275979 166461 275980
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 161979 238644 162045 238645
rect 161979 238580 161980 238644
rect 162044 238580 162045 238644
rect 161979 238579 162045 238580
rect 163794 237454 164414 272898
rect 166211 243540 166277 243541
rect 166211 243476 166212 243540
rect 166276 243476 166277 243540
rect 166211 243475 166277 243476
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 160691 180028 160757 180029
rect 160691 179964 160692 180028
rect 160756 179964 160757 180028
rect 160691 179963 160757 179964
rect 163794 176600 164414 200898
rect 166214 180165 166274 243475
rect 166398 220829 166458 275979
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 166395 220828 166461 220829
rect 166395 220764 166396 220828
rect 166460 220764 166461 220828
rect 166395 220763 166461 220764
rect 168294 205954 168914 241398
rect 169710 231845 169770 295563
rect 171731 265572 171797 265573
rect 171731 265508 171732 265572
rect 171796 265508 171797 265572
rect 171731 265507 171797 265508
rect 169707 231844 169773 231845
rect 169707 231780 169708 231844
rect 169772 231780 169773 231844
rect 169707 231779 169773 231780
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 166395 182204 166461 182205
rect 166395 182140 166396 182204
rect 166460 182140 166461 182204
rect 166395 182139 166461 182140
rect 166211 180164 166277 180165
rect 166211 180100 166212 180164
rect 166276 180100 166277 180164
rect 166211 180099 166277 180100
rect 166211 178124 166277 178125
rect 166211 178060 166212 178124
rect 166276 178060 166277 178124
rect 166211 178059 166277 178060
rect 135670 175070 135780 175130
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 166214 154597 166274 178059
rect 166398 163165 166458 182139
rect 167683 178260 167749 178261
rect 167683 178196 167684 178260
rect 167748 178196 167749 178260
rect 167683 178195 167749 178196
rect 167499 176900 167565 176901
rect 167499 176836 167500 176900
rect 167564 176836 167565 176900
rect 167499 176835 167565 176836
rect 166395 163164 166461 163165
rect 166395 163100 166396 163164
rect 166460 163100 166461 163164
rect 166395 163099 166461 163100
rect 167502 157453 167562 176835
rect 167686 161533 167746 178195
rect 168294 169954 168914 205398
rect 169707 181660 169773 181661
rect 169707 181596 169708 181660
rect 169772 181596 169773 181660
rect 169707 181595 169773 181596
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 167683 161532 167749 161533
rect 167683 161468 167684 161532
rect 167748 161468 167749 161532
rect 167683 161467 167749 161468
rect 167499 157452 167565 157453
rect 167499 157388 167500 157452
rect 167564 157388 167565 157452
rect 167499 157387 167565 157388
rect 166211 154596 166277 154597
rect 166211 154532 166212 154596
rect 166276 154532 166277 154596
rect 166211 154531 166277 154532
rect 69072 151954 69420 151986
rect 69072 151718 69128 151954
rect 69364 151718 69420 151954
rect 69072 151634 69420 151718
rect 69072 151398 69128 151634
rect 69364 151398 69420 151634
rect 69072 151366 69420 151398
rect 164136 151954 164484 151986
rect 164136 151718 164192 151954
rect 164428 151718 164484 151954
rect 164136 151634 164484 151718
rect 164136 151398 164192 151634
rect 164428 151398 164484 151634
rect 164136 151366 164484 151398
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 167499 143716 167565 143717
rect 167499 143652 167500 143716
rect 167564 143652 167565 143716
rect 167499 143651 167565 143652
rect 166211 131204 166277 131205
rect 166211 131140 166212 131204
rect 166276 131140 166277 131204
rect 166211 131139 166277 131140
rect 69072 115954 69420 115986
rect 69072 115718 69128 115954
rect 69364 115718 69420 115954
rect 69072 115634 69420 115718
rect 69072 115398 69128 115634
rect 69364 115398 69420 115634
rect 69072 115366 69420 115398
rect 164136 115954 164484 115986
rect 164136 115718 164192 115954
rect 164428 115718 164484 115954
rect 164136 115634 164484 115718
rect 164136 115398 164192 115634
rect 164428 115398 164484 115634
rect 164136 115366 164484 115398
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85682 94890
rect 86624 94830 86786 94890
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 70954 69914 93100
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 75454 74414 93100
rect 74766 92445 74826 94830
rect 74763 92444 74829 92445
rect 74763 92380 74764 92444
rect 74828 92380 74829 92444
rect 74763 92379 74829 92380
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 79954 78914 93100
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 84454 83414 93100
rect 84334 91221 84394 94830
rect 85622 92445 85682 94830
rect 85619 92444 85685 92445
rect 85619 92380 85620 92444
rect 85684 92380 85685 92444
rect 85619 92379 85685 92380
rect 86726 91221 86786 94830
rect 87094 94830 88044 94890
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 87094 91221 87154 94830
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 87091 91220 87157 91221
rect 87091 91156 87092 91220
rect 87156 91156 87157 91220
rect 87091 91155 87157 91156
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 88954 87914 93100
rect 88934 91765 88994 94830
rect 88931 91764 88997 91765
rect 88931 91700 88932 91764
rect 88996 91700 88997 91764
rect 88931 91699 88997 91700
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96170 94890
rect 96688 94830 96906 94890
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 99136 94830 99298 94890
rect 99544 94830 99666 94890
rect 91326 91221 91386 94830
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 92445 93962 94830
rect 93899 92444 93965 92445
rect 93899 92380 93900 92444
rect 93964 92380 93965 92444
rect 93899 92379 93965 92380
rect 95006 91221 95066 94830
rect 96110 91221 96170 94830
rect 96846 93870 96906 94830
rect 96846 93810 97090 93870
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 96107 91220 96173 91221
rect 96107 91156 96108 91220
rect 96172 91156 96173 91220
rect 96107 91155 96173 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 61954 96914 93100
rect 97030 91357 97090 93810
rect 97027 91356 97093 91357
rect 97027 91292 97028 91356
rect 97092 91292 97093 91356
rect 97027 91291 97093 91292
rect 97214 91221 97274 94830
rect 98134 91357 98194 94830
rect 98502 91493 98562 94830
rect 98499 91492 98565 91493
rect 98499 91428 98500 91492
rect 98564 91428 98565 91492
rect 98499 91427 98565 91428
rect 98131 91356 98197 91357
rect 98131 91292 98132 91356
rect 98196 91292 98197 91356
rect 98131 91291 98197 91292
rect 99238 91221 99298 94830
rect 99606 91221 99666 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 101690 94890
rect 100526 91221 100586 94830
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 99235 91220 99301 91221
rect 99235 91156 99236 91220
rect 99300 91156 99301 91220
rect 99235 91155 99301 91156
rect 99603 91220 99669 91221
rect 99603 91156 99604 91220
rect 99668 91156 99669 91220
rect 99603 91155 99669 91156
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 66454 101414 93100
rect 101630 91221 101690 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 92445 101874 94830
rect 101998 93533 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 101995 93532 102061 93533
rect 101995 93468 101996 93532
rect 102060 93468 102061 93532
rect 101995 93467 102061 93468
rect 101811 92444 101877 92445
rect 101811 92380 101812 92444
rect 101876 92380 101877 92444
rect 101811 92379 101877 92380
rect 102918 91221 102978 94830
rect 103286 91221 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 104440 94830 104634 94890
rect 104206 91629 104266 94830
rect 104203 91628 104269 91629
rect 104203 91564 104204 91628
rect 104268 91564 104269 91628
rect 104203 91563 104269 91564
rect 104574 91221 104634 94830
rect 105126 94830 105452 94890
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 105664 94830 106106 94890
rect 105126 91221 105186 94830
rect 101627 91220 101693 91221
rect 101627 91156 101628 91220
rect 101692 91156 101693 91220
rect 101627 91155 101693 91156
rect 102915 91220 102981 91221
rect 102915 91156 102916 91220
rect 102980 91156 102981 91220
rect 102915 91155 102981 91156
rect 103283 91220 103349 91221
rect 103283 91156 103284 91220
rect 103348 91156 103349 91220
rect 103283 91155 103349 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105123 91220 105189 91221
rect 105123 91156 105124 91220
rect 105188 91156 105189 91220
rect 105123 91155 105189 91156
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 70954 105914 93100
rect 106046 92173 106106 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 106043 92172 106109 92173
rect 106043 92108 106044 92172
rect 106108 92108 106109 92172
rect 106043 92107 106109 92108
rect 106414 91221 106474 94830
rect 106782 91629 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 107702 93533 107762 94830
rect 108070 93805 108130 94830
rect 109064 94757 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109472 94830 109602 94890
rect 109061 94756 109127 94757
rect 109061 94692 109062 94756
rect 109126 94692 109127 94756
rect 109061 94691 109127 94692
rect 108067 93804 108133 93805
rect 108067 93740 108068 93804
rect 108132 93740 108133 93804
rect 108067 93739 108133 93740
rect 107699 93532 107765 93533
rect 107699 93468 107700 93532
rect 107764 93468 107765 93532
rect 107699 93467 107765 93468
rect 106779 91628 106845 91629
rect 106779 91564 106780 91628
rect 106844 91564 106845 91628
rect 106779 91563 106845 91564
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 106411 91220 106477 91221
rect 106411 91156 106412 91220
rect 106476 91156 106477 91220
rect 106411 91155 106477 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 91221 111258 94830
rect 111934 92309 111994 94830
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113144 94830 113282 94890
rect 111931 92308 111997 92309
rect 111931 92244 111932 92308
rect 111996 92244 111997 92308
rect 111931 92243 111997 92244
rect 112302 91765 112362 94830
rect 112299 91764 112365 91765
rect 112299 91700 112300 91764
rect 112364 91700 112365 91764
rect 112299 91699 112365 91700
rect 113222 91221 113282 94830
rect 113688 94757 113748 95200
rect 114368 94890 114428 95200
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 115122 94890
rect 113685 94756 113751 94757
rect 113685 94692 113686 94756
rect 113750 94692 113751 94756
rect 113685 94691 113751 94692
rect 114326 93941 114386 94830
rect 114323 93940 114389 93941
rect 114323 93876 114324 93940
rect 114388 93876 114389 93940
rect 114323 93875 114389 93876
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 113219 91220 113285 91221
rect 113219 91156 113220 91220
rect 113284 91156 113285 91220
rect 113219 91155 113285 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 79954 114914 93100
rect 115062 92445 115122 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 92445 115490 94830
rect 115059 92444 115125 92445
rect 115059 92380 115060 92444
rect 115124 92380 115125 92444
rect 115059 92379 115125 92380
rect 115427 92444 115493 92445
rect 115427 92380 115428 92444
rect 115492 92380 115493 92444
rect 115427 92379 115493 92380
rect 115798 91221 115858 94830
rect 116718 91221 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 117086 91221 117146 94830
rect 118006 91221 118066 94830
rect 118190 91357 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119294 93261 119354 94830
rect 119291 93260 119357 93261
rect 119291 93196 119292 93260
rect 119356 93196 119357 93260
rect 119291 93195 119357 93196
rect 118187 91356 118253 91357
rect 118187 91292 118188 91356
rect 118252 91292 118253 91356
rect 118187 91291 118253 91292
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 116715 91220 116781 91221
rect 116715 91156 116716 91220
rect 116780 91156 116781 91220
rect 116715 91155 116781 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 118003 91220 118069 91221
rect 118003 91156 118004 91220
rect 118068 91156 118069 91220
rect 118003 91155 118069 91156
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 84454 119414 93100
rect 119662 91221 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 121984 94830 122114 94890
rect 120214 92445 120274 94830
rect 120211 92444 120277 92445
rect 120211 92380 120212 92444
rect 120276 92380 120277 92444
rect 120211 92379 120277 92380
rect 120582 91221 120642 94830
rect 121686 93669 121746 94830
rect 121683 93668 121749 93669
rect 121683 93604 121684 93668
rect 121748 93604 121749 93668
rect 121683 93603 121749 93604
rect 122054 91221 122114 94830
rect 122800 93870 122860 95200
rect 123208 94890 123268 95200
rect 122606 93810 122860 93870
rect 122974 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 122974 91765 123034 94830
rect 122971 91764 123037 91765
rect 122971 91700 122972 91764
rect 123036 91700 123037 91764
rect 122971 91699 123037 91700
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 119659 91220 119725 91221
rect 119659 91156 119660 91220
rect 119724 91156 119725 91220
rect 119659 91155 119725 91156
rect 120579 91220 120645 91221
rect 120579 91156 120580 91220
rect 120644 91156 120645 91220
rect 120579 91155 120645 91156
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 88954 123914 93100
rect 124078 92445 124138 94830
rect 124446 93533 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125978 94890
rect 124443 93532 124509 93533
rect 124443 93468 124444 93532
rect 124508 93468 124509 93532
rect 124443 93467 124509 93468
rect 124075 92444 124141 92445
rect 124075 92380 124076 92444
rect 124140 92380 124141 92444
rect 124075 92379 124141 92380
rect 125366 91221 125426 94830
rect 125918 92445 125978 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125915 92444 125981 92445
rect 125915 92380 125916 92444
rect 125980 92380 125981 92444
rect 125915 92379 125981 92380
rect 126470 91629 126530 94830
rect 126467 91628 126533 91629
rect 126467 91564 126468 91628
rect 126532 91564 126533 91628
rect 126467 91563 126533 91564
rect 126654 91221 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 127574 91221 127634 94830
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 91221 130762 94830
rect 131912 94757 131972 95200
rect 133136 94890 133196 95200
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 135730 94890
rect 131909 94756 131975 94757
rect 131909 94692 131910 94756
rect 131974 94692 131975 94756
rect 131909 94691 131975 94692
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 93100
rect 133094 92445 133154 94830
rect 133091 92444 133157 92445
rect 133091 92380 133092 92444
rect 133156 92380 133157 92444
rect 133091 92379 133157 92380
rect 134382 91221 134442 94830
rect 135670 91221 135730 94830
rect 151310 94830 151556 94890
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 135667 91220 135733 91221
rect 135667 91156 135668 91220
rect 135732 91156 135733 91220
rect 135667 91155 135733 91156
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 93100
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 70954 141914 93100
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 79954 150914 93100
rect 151310 91765 151370 94830
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151904 94757 151964 95200
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151765 94691 151831 94692
rect 151901 94756 151967 94757
rect 151901 94692 151902 94756
rect 151966 94692 151967 94756
rect 151901 94691 151967 94692
rect 151632 94150 151738 94210
rect 151678 92445 151738 94150
rect 151675 92444 151741 92445
rect 151675 92380 151676 92444
rect 151740 92380 151741 92444
rect 151675 92379 151741 92380
rect 151307 91764 151373 91765
rect 151307 91700 151308 91764
rect 151372 91700 151373 91764
rect 151307 91699 151373 91700
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 84454 155414 93100
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 88954 159914 93100
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 93100
rect 166214 86869 166274 131139
rect 166395 97204 166461 97205
rect 166395 97140 166396 97204
rect 166460 97140 166461 97204
rect 166395 97139 166461 97140
rect 166398 92309 166458 97139
rect 166395 92308 166461 92309
rect 166395 92244 166396 92308
rect 166460 92244 166461 92308
rect 166395 92243 166461 92244
rect 167502 91085 167562 143651
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 167683 132836 167749 132837
rect 167683 132772 167684 132836
rect 167748 132772 167749 132836
rect 167683 132771 167749 132772
rect 167686 93805 167746 132771
rect 168294 97954 168914 133398
rect 169155 128620 169221 128621
rect 169155 128556 169156 128620
rect 169220 128556 169221 128620
rect 169155 128555 169221 128556
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 167683 93804 167749 93805
rect 167683 93740 167684 93804
rect 167748 93740 167749 93804
rect 167683 93739 167749 93740
rect 167499 91084 167565 91085
rect 167499 91020 167500 91084
rect 167564 91020 167565 91084
rect 167499 91019 167565 91020
rect 166211 86868 166277 86869
rect 166211 86804 166212 86868
rect 166276 86804 166277 86868
rect 166211 86803 166277 86804
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 97398
rect 169158 78573 169218 128555
rect 169155 78572 169221 78573
rect 169155 78508 169156 78572
rect 169220 78508 169221 78572
rect 169155 78507 169221 78508
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 169710 3365 169770 181595
rect 170259 133924 170325 133925
rect 170259 133860 170260 133924
rect 170324 133860 170325 133924
rect 170259 133859 170325 133860
rect 170262 84149 170322 133859
rect 171734 95981 171794 265507
rect 172286 255237 172346 359347
rect 172794 354454 173414 389898
rect 177294 394954 177914 403000
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 181794 399454 182414 403000
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 180011 390012 180077 390013
rect 180011 389948 180012 390012
rect 180076 389948 180077 390012
rect 180011 389947 180077 389948
rect 178539 387020 178605 387021
rect 178539 386956 178540 387020
rect 178604 386956 178605 387020
rect 178539 386955 178605 386956
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177067 355332 177133 355333
rect 177067 355268 177068 355332
rect 177132 355268 177133 355332
rect 177067 355267 177133 355268
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 176515 350164 176581 350165
rect 176515 350100 176516 350164
rect 176580 350100 176581 350164
rect 176515 350099 176581 350100
rect 176331 339284 176397 339285
rect 176331 339220 176332 339284
rect 176396 339220 176397 339284
rect 176331 339219 176397 339220
rect 175043 321604 175109 321605
rect 175043 321540 175044 321604
rect 175108 321540 175109 321604
rect 175043 321539 175109 321540
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 173571 294540 173637 294541
rect 173571 294476 173572 294540
rect 173636 294476 173637 294540
rect 173571 294475 173637 294476
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172283 255236 172349 255237
rect 172283 255172 172284 255236
rect 172348 255172 172349 255236
rect 172283 255171 172349 255172
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 171731 95980 171797 95981
rect 171731 95916 171732 95980
rect 171796 95916 171797 95980
rect 171731 95915 171797 95916
rect 170259 84148 170325 84149
rect 170259 84084 170260 84148
rect 170324 84084 170325 84148
rect 170259 84083 170325 84084
rect 172794 66454 173414 101898
rect 173574 93805 173634 294475
rect 174491 293996 174557 293997
rect 174491 293932 174492 293996
rect 174556 293932 174557 293996
rect 174491 293931 174557 293932
rect 173571 93804 173637 93805
rect 173571 93740 173572 93804
rect 173636 93740 173637 93804
rect 173571 93739 173637 93740
rect 174494 92445 174554 293931
rect 174491 92444 174557 92445
rect 174491 92380 174492 92444
rect 174556 92380 174557 92444
rect 174491 92379 174557 92380
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 169707 3364 169773 3365
rect 169707 3300 169708 3364
rect 169772 3300 169773 3364
rect 169707 3299 169773 3300
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 175046 6221 175106 321539
rect 176334 39269 176394 339219
rect 176331 39268 176397 39269
rect 176331 39204 176332 39268
rect 176396 39204 176397 39268
rect 176331 39203 176397 39204
rect 175043 6220 175109 6221
rect 175043 6156 175044 6220
rect 175108 6156 175109 6220
rect 175043 6155 175109 6156
rect 176518 2005 176578 350099
rect 177070 262173 177130 355267
rect 177294 322954 177914 358398
rect 178542 349757 178602 386955
rect 179827 352612 179893 352613
rect 179827 352548 179828 352612
rect 179892 352610 179893 352612
rect 180014 352610 180074 389947
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 357154 182414 362898
rect 213294 394954 213914 403000
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 357154 213914 358398
rect 217794 399454 218414 403000
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 242942 380221 243002 567150
rect 244227 553348 244293 553349
rect 244227 553284 244228 553348
rect 244292 553284 244293 553348
rect 244227 553283 244293 553284
rect 243307 407284 243373 407285
rect 243307 407220 243308 407284
rect 243372 407220 243373 407284
rect 243307 407219 243373 407220
rect 243310 403613 243370 407219
rect 243307 403612 243373 403613
rect 243307 403548 243308 403612
rect 243372 403548 243373 403612
rect 243307 403547 243373 403548
rect 244230 389877 244290 553283
rect 244411 546548 244477 546549
rect 244411 546484 244412 546548
rect 244476 546484 244477 546548
rect 244411 546483 244477 546484
rect 244414 400893 244474 546483
rect 245699 529548 245765 529549
rect 245699 529484 245700 529548
rect 245764 529484 245765 529548
rect 245699 529483 245765 529484
rect 244411 400892 244477 400893
rect 244411 400828 244412 400892
rect 244476 400828 244477 400892
rect 244411 400827 244477 400828
rect 244227 389876 244293 389877
rect 244227 389812 244228 389876
rect 244292 389812 244293 389876
rect 244227 389811 244293 389812
rect 242939 380220 243005 380221
rect 242939 380156 242940 380220
rect 243004 380156 243005 380220
rect 242939 380155 243005 380156
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 357154 218414 362898
rect 245702 362269 245762 529483
rect 245883 489428 245949 489429
rect 245883 489364 245884 489428
rect 245948 489364 245949 489428
rect 245883 489363 245949 489364
rect 245886 401029 245946 489363
rect 245883 401028 245949 401029
rect 245883 400964 245884 401028
rect 245948 400964 245949 401028
rect 245883 400963 245949 400964
rect 246990 380357 247050 569603
rect 247174 405517 247234 585379
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 247171 405516 247237 405517
rect 247171 405452 247172 405516
rect 247236 405452 247237 405516
rect 247171 405451 247237 405452
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 246987 380356 247053 380357
rect 246987 380292 246988 380356
rect 247052 380292 247053 380356
rect 246987 380291 247053 380292
rect 245699 362268 245765 362269
rect 245699 362204 245700 362268
rect 245764 362204 245765 362268
rect 245699 362203 245765 362204
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 357154 249914 358398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 357154 254414 362898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 357154 258914 367398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 357154 263414 371898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 357154 267914 376398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 357154 272414 380898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 357154 276914 385398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 357154 281414 389898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 357154 285914 358398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 357154 290414 362898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 295379 578916 295445 578917
rect 295379 578852 295380 578916
rect 295444 578852 295445 578916
rect 295379 578851 295445 578852
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 295011 375324 295077 375325
rect 295011 375260 295012 375324
rect 295076 375260 295077 375324
rect 295011 375259 295077 375260
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 293907 357372 293973 357373
rect 293907 357308 293908 357372
rect 293972 357308 293973 357372
rect 293907 357307 293973 357308
rect 292619 356148 292685 356149
rect 292619 356084 292620 356148
rect 292684 356084 292685 356148
rect 292619 356083 292685 356084
rect 179892 352550 180074 352610
rect 179892 352548 179893 352550
rect 179827 352547 179893 352548
rect 178539 349756 178605 349757
rect 178539 349692 178540 349756
rect 178604 349692 178605 349756
rect 178539 349691 178605 349692
rect 199568 331954 199888 331986
rect 199568 331718 199610 331954
rect 199846 331718 199888 331954
rect 199568 331634 199888 331718
rect 199568 331398 199610 331634
rect 199846 331398 199888 331634
rect 199568 331366 199888 331398
rect 230288 331954 230608 331986
rect 230288 331718 230330 331954
rect 230566 331718 230608 331954
rect 230288 331634 230608 331718
rect 230288 331398 230330 331634
rect 230566 331398 230608 331634
rect 230288 331366 230608 331398
rect 261008 331954 261328 331986
rect 261008 331718 261050 331954
rect 261286 331718 261328 331954
rect 261008 331634 261328 331718
rect 261008 331398 261050 331634
rect 261286 331398 261328 331634
rect 261008 331366 261328 331398
rect 179275 327724 179341 327725
rect 179275 327660 179276 327724
rect 179340 327660 179341 327724
rect 179275 327659 179341 327660
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177067 262172 177133 262173
rect 177067 262108 177068 262172
rect 177132 262108 177133 262172
rect 177067 262107 177133 262108
rect 177067 259724 177133 259725
rect 177067 259660 177068 259724
rect 177132 259660 177133 259724
rect 177067 259659 177133 259660
rect 177070 50285 177130 259659
rect 177294 250954 177914 286398
rect 179091 279580 179157 279581
rect 179091 279516 179092 279580
rect 179156 279516 179157 279580
rect 179091 279515 179157 279516
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 179094 226949 179154 279515
rect 179278 256733 179338 327659
rect 184208 327454 184528 327486
rect 184208 327218 184250 327454
rect 184486 327218 184528 327454
rect 184208 327134 184528 327218
rect 184208 326898 184250 327134
rect 184486 326898 184528 327134
rect 184208 326866 184528 326898
rect 214928 327454 215248 327486
rect 214928 327218 214970 327454
rect 215206 327218 215248 327454
rect 214928 327134 215248 327218
rect 214928 326898 214970 327134
rect 215206 326898 215248 327134
rect 214928 326866 215248 326898
rect 245648 327454 245968 327486
rect 245648 327218 245690 327454
rect 245926 327218 245968 327454
rect 245648 327134 245968 327218
rect 245648 326898 245690 327134
rect 245926 326898 245968 327134
rect 245648 326866 245968 326898
rect 276368 327454 276688 327486
rect 276368 327218 276410 327454
rect 276646 327218 276688 327454
rect 276368 327134 276688 327218
rect 276368 326898 276410 327134
rect 276646 326898 276688 327134
rect 276368 326866 276688 326898
rect 292622 303517 292682 356083
rect 293171 309092 293237 309093
rect 293171 309028 293172 309092
rect 293236 309028 293237 309092
rect 293171 309027 293237 309028
rect 292619 303516 292685 303517
rect 292619 303452 292620 303516
rect 292684 303452 292685 303516
rect 292619 303451 292685 303452
rect 199568 295954 199888 295986
rect 199568 295718 199610 295954
rect 199846 295718 199888 295954
rect 199568 295634 199888 295718
rect 199568 295398 199610 295634
rect 199846 295398 199888 295634
rect 199568 295366 199888 295398
rect 230288 295954 230608 295986
rect 230288 295718 230330 295954
rect 230566 295718 230608 295954
rect 230288 295634 230608 295718
rect 230288 295398 230330 295634
rect 230566 295398 230608 295634
rect 230288 295366 230608 295398
rect 261008 295954 261328 295986
rect 261008 295718 261050 295954
rect 261286 295718 261328 295954
rect 261008 295634 261328 295718
rect 261008 295398 261050 295634
rect 261286 295398 261328 295634
rect 261008 295366 261328 295398
rect 184208 291454 184528 291486
rect 184208 291218 184250 291454
rect 184486 291218 184528 291454
rect 184208 291134 184528 291218
rect 184208 290898 184250 291134
rect 184486 290898 184528 291134
rect 184208 290866 184528 290898
rect 214928 291454 215248 291486
rect 214928 291218 214970 291454
rect 215206 291218 215248 291454
rect 214928 291134 215248 291218
rect 214928 290898 214970 291134
rect 215206 290898 215248 291134
rect 214928 290866 215248 290898
rect 245648 291454 245968 291486
rect 245648 291218 245690 291454
rect 245926 291218 245968 291454
rect 245648 291134 245968 291218
rect 245648 290898 245690 291134
rect 245926 290898 245968 291134
rect 245648 290866 245968 290898
rect 276368 291454 276688 291486
rect 276368 291218 276410 291454
rect 276646 291218 276688 291454
rect 276368 291134 276688 291218
rect 276368 290898 276410 291134
rect 276646 290898 276688 291134
rect 276368 290866 276688 290898
rect 292619 281756 292685 281757
rect 292619 281692 292620 281756
rect 292684 281692 292685 281756
rect 292619 281691 292685 281692
rect 199568 259954 199888 259986
rect 199568 259718 199610 259954
rect 199846 259718 199888 259954
rect 199568 259634 199888 259718
rect 199568 259398 199610 259634
rect 199846 259398 199888 259634
rect 199568 259366 199888 259398
rect 230288 259954 230608 259986
rect 230288 259718 230330 259954
rect 230566 259718 230608 259954
rect 230288 259634 230608 259718
rect 230288 259398 230330 259634
rect 230566 259398 230608 259634
rect 230288 259366 230608 259398
rect 261008 259954 261328 259986
rect 261008 259718 261050 259954
rect 261286 259718 261328 259954
rect 261008 259634 261328 259718
rect 261008 259398 261050 259634
rect 261286 259398 261328 259634
rect 261008 259366 261328 259398
rect 179275 256732 179341 256733
rect 179275 256668 179276 256732
rect 179340 256668 179341 256732
rect 179275 256667 179341 256668
rect 184208 255454 184528 255486
rect 184208 255218 184250 255454
rect 184486 255218 184528 255454
rect 184208 255134 184528 255218
rect 184208 254898 184250 255134
rect 184486 254898 184528 255134
rect 184208 254866 184528 254898
rect 214928 255454 215248 255486
rect 214928 255218 214970 255454
rect 215206 255218 215248 255454
rect 214928 255134 215248 255218
rect 214928 254898 214970 255134
rect 215206 254898 215248 255134
rect 214928 254866 215248 254898
rect 245648 255454 245968 255486
rect 245648 255218 245690 255454
rect 245926 255218 245968 255454
rect 245648 255134 245968 255218
rect 245648 254898 245690 255134
rect 245926 254898 245968 255134
rect 245648 254866 245968 254898
rect 276368 255454 276688 255486
rect 276368 255218 276410 255454
rect 276646 255218 276688 255454
rect 276368 255134 276688 255218
rect 276368 254898 276410 255134
rect 276646 254898 276688 255134
rect 276368 254866 276688 254898
rect 179275 248164 179341 248165
rect 179275 248100 179276 248164
rect 179340 248100 179341 248164
rect 179275 248099 179341 248100
rect 179091 226948 179157 226949
rect 179091 226884 179092 226948
rect 179156 226884 179157 226948
rect 179091 226883 179157 226884
rect 178907 226404 178973 226405
rect 178907 226340 178908 226404
rect 178972 226340 178973 226404
rect 178907 226339 178973 226340
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 178910 89045 178970 226339
rect 178907 89044 178973 89045
rect 178907 88980 178908 89044
rect 178972 88980 178973 89044
rect 178907 88979 178973 88980
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177067 50284 177133 50285
rect 177067 50220 177068 50284
rect 177132 50220 177133 50284
rect 177067 50219 177133 50220
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 176515 2004 176581 2005
rect 176515 1940 176516 2004
rect 176580 1940 176581 2004
rect 176515 1939 176581 1940
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 -7066 177914 34398
rect 179278 21317 179338 248099
rect 179643 243676 179709 243677
rect 179643 243612 179644 243676
rect 179708 243612 179709 243676
rect 179643 243611 179709 243612
rect 179646 79389 179706 243611
rect 179827 243540 179893 243541
rect 179827 243476 179828 243540
rect 179892 243476 179893 243540
rect 179827 243475 179893 243476
rect 179830 231845 179890 243475
rect 292622 239189 292682 281691
rect 292619 239188 292685 239189
rect 292619 239124 292620 239188
rect 292684 239124 292685 239188
rect 292619 239123 292685 239124
rect 179827 231844 179893 231845
rect 179827 231780 179828 231844
rect 179892 231780 179893 231844
rect 179827 231779 179893 231780
rect 181794 219454 182414 238000
rect 184795 237420 184861 237421
rect 184795 237356 184796 237420
rect 184860 237356 184861 237420
rect 184795 237355 184861 237356
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 179643 79388 179709 79389
rect 179643 79324 179644 79388
rect 179708 79324 179709 79388
rect 179643 79323 179709 79324
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 179275 21316 179341 21317
rect 179275 21252 179276 21316
rect 179340 21252 179341 21316
rect 179275 21251 179341 21252
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 3454 182414 38898
rect 184798 18733 184858 237355
rect 186294 223954 186914 238000
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 184795 18732 184861 18733
rect 184795 18668 184796 18732
rect 184860 18668 184861 18732
rect 184795 18667 184861 18668
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228454 191414 238000
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 232954 195914 238000
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 237454 200414 238000
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 238000
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 238000
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 238000
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 217794 219454 218414 238000
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 222294 223954 222914 238000
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 178000 222914 187398
rect 226794 228454 227414 238000
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 178000 227414 191898
rect 231294 232954 231914 238000
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 178000 231914 196398
rect 235794 237454 236414 238000
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 249294 214954 249914 238000
rect 252507 222868 252573 222869
rect 252507 222804 252508 222868
rect 252572 222804 252573 222868
rect 252507 222803 252573 222804
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249011 178940 249077 178941
rect 249011 178876 249012 178940
rect 249076 178876 249077 178940
rect 249011 178875 249077 178876
rect 249014 177850 249074 178875
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 178000 249914 178398
rect 249014 177790 249442 177850
rect 249195 177580 249261 177581
rect 249195 177516 249196 177580
rect 249260 177516 249261 177580
rect 249195 177515 249261 177516
rect 249198 174317 249258 177515
rect 249195 174316 249261 174317
rect 249195 174252 249196 174316
rect 249260 174252 249261 174316
rect 249195 174251 249261 174252
rect 249382 173365 249442 177790
rect 249379 173364 249445 173365
rect 249379 173300 249380 173364
rect 249444 173300 249445 173364
rect 249379 173299 249445 173300
rect 252510 155413 252570 222803
rect 253794 219454 254414 238000
rect 256739 225588 256805 225589
rect 256739 225524 256740 225588
rect 256804 225524 256805 225588
rect 256739 225523 256805 225524
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 255451 186420 255517 186421
rect 255451 186356 255452 186420
rect 255516 186356 255517 186420
rect 255451 186355 255517 186356
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 252507 155412 252573 155413
rect 252507 155348 252508 155412
rect 252572 155348 252573 155412
rect 252507 155347 252573 155348
rect 227874 151954 228194 151986
rect 227874 151718 227916 151954
rect 228152 151718 228194 151954
rect 227874 151634 228194 151718
rect 227874 151398 227916 151634
rect 228152 151398 228194 151634
rect 227874 151366 228194 151398
rect 237805 151954 238125 151986
rect 237805 151718 237847 151954
rect 238083 151718 238125 151954
rect 237805 151634 238125 151718
rect 237805 151398 237847 151634
rect 238083 151398 238125 151634
rect 237805 151366 238125 151398
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 253794 147454 254414 182898
rect 255267 181524 255333 181525
rect 255267 181460 255268 181524
rect 255332 181460 255333 181524
rect 255267 181459 255333 181460
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 251771 141132 251837 141133
rect 251771 141068 251772 141132
rect 251836 141068 251837 141132
rect 251771 141067 251837 141068
rect 227874 115954 228194 115986
rect 227874 115718 227916 115954
rect 228152 115718 228194 115954
rect 227874 115634 228194 115718
rect 227874 115398 227916 115634
rect 228152 115398 228194 115634
rect 227874 115366 228194 115398
rect 237805 115954 238125 115986
rect 237805 115718 237847 115954
rect 238083 115718 238125 115954
rect 237805 115634 238125 115718
rect 237805 115398 237847 115634
rect 238083 115398 238125 115634
rect 237805 115366 238125 115398
rect 251774 113117 251834 141067
rect 251955 115156 252021 115157
rect 251955 115092 251956 115156
rect 252020 115092 252021 115156
rect 251955 115091 252021 115092
rect 251771 113116 251837 113117
rect 251771 113052 251772 113116
rect 251836 113052 251837 113116
rect 251771 113051 251837 113052
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 242771 110866 243091 110898
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 251958 98021 252018 115091
rect 253794 111454 254414 146898
rect 255270 139909 255330 181459
rect 255454 147933 255514 186355
rect 256742 169829 256802 225523
rect 258294 223954 258914 238000
rect 262794 228454 263414 238000
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 259499 224228 259565 224229
rect 259499 224164 259500 224228
rect 259564 224164 259565 224228
rect 259499 224163 259565 224164
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 257843 194036 257909 194037
rect 257843 193972 257844 194036
rect 257908 193972 257909 194036
rect 257843 193971 257909 193972
rect 256923 178668 256989 178669
rect 256923 178604 256924 178668
rect 256988 178604 256989 178668
rect 256923 178603 256989 178604
rect 256739 169828 256805 169829
rect 256739 169764 256740 169828
rect 256804 169764 256805 169828
rect 256739 169763 256805 169764
rect 256926 164253 256986 178603
rect 256923 164252 256989 164253
rect 256923 164188 256924 164252
rect 256988 164188 256989 164252
rect 256923 164187 256989 164188
rect 255451 147932 255517 147933
rect 255451 147868 255452 147932
rect 255516 147868 255517 147932
rect 255451 147867 255517 147868
rect 257846 146301 257906 193971
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 257843 146300 257909 146301
rect 257843 146236 257844 146300
rect 257908 146236 257909 146300
rect 257843 146235 257909 146236
rect 255267 139908 255333 139909
rect 255267 139844 255268 139908
rect 255332 139844 255333 139908
rect 255267 139843 255333 139844
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 251955 98020 252021 98021
rect 251955 97956 251956 98020
rect 252020 97956 252021 98020
rect 251955 97955 252021 97956
rect 250115 97068 250181 97069
rect 250115 97004 250116 97068
rect 250180 97004 250181 97068
rect 250115 97003 250181 97004
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 79954 222914 94000
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 84454 227414 94000
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 88954 231914 94000
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 61954 240914 94000
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 66454 245414 94000
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 70954 249914 94000
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 250118 16557 250178 97003
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 250115 16556 250181 16557
rect 250115 16492 250116 16556
rect 250180 16492 250181 16556
rect 250115 16491 250181 16492
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 115954 258914 151398
rect 259502 138957 259562 224163
rect 260971 202332 261037 202333
rect 260971 202268 260972 202332
rect 261036 202268 261037 202332
rect 260971 202267 261037 202268
rect 260787 191044 260853 191045
rect 260787 190980 260788 191044
rect 260852 190980 260853 191044
rect 260787 190979 260853 190980
rect 259683 178804 259749 178805
rect 259683 178740 259684 178804
rect 259748 178740 259749 178804
rect 259683 178739 259749 178740
rect 259686 141269 259746 178739
rect 260790 171150 260850 190979
rect 260974 173909 261034 202267
rect 262794 192454 263414 227898
rect 267294 232954 267914 238000
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 265019 204916 265085 204917
rect 265019 204852 265020 204916
rect 265084 204852 265085 204916
rect 265019 204851 265085 204852
rect 263731 192540 263797 192541
rect 263731 192476 263732 192540
rect 263796 192476 263797 192540
rect 263731 192475 263797 192476
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262259 176084 262325 176085
rect 262259 176020 262260 176084
rect 262324 176020 262325 176084
rect 262259 176019 262325 176020
rect 260971 173908 261037 173909
rect 260971 173844 260972 173908
rect 261036 173844 261037 173908
rect 260971 173843 261037 173844
rect 261339 171460 261405 171461
rect 261339 171396 261340 171460
rect 261404 171396 261405 171460
rect 261339 171395 261405 171396
rect 260790 171090 261034 171150
rect 260974 142765 261034 171090
rect 260971 142764 261037 142765
rect 260971 142700 260972 142764
rect 261036 142700 261037 142764
rect 260971 142699 261037 142700
rect 261342 141541 261402 171395
rect 262262 157861 262322 176019
rect 262259 157860 262325 157861
rect 262259 157796 262260 157860
rect 262324 157796 262325 157860
rect 262259 157795 262325 157796
rect 262794 156454 263414 191898
rect 263547 188460 263613 188461
rect 263547 188396 263548 188460
rect 263612 188396 263613 188460
rect 263547 188395 263613 188396
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 261339 141540 261405 141541
rect 261339 141476 261340 141540
rect 261404 141476 261405 141540
rect 261339 141475 261405 141476
rect 259683 141268 259749 141269
rect 259683 141204 259684 141268
rect 259748 141204 259749 141268
rect 259683 141203 259749 141204
rect 261339 139772 261405 139773
rect 261339 139708 261340 139772
rect 261404 139708 261405 139772
rect 261339 139707 261405 139708
rect 259499 138956 259565 138957
rect 259499 138892 259500 138956
rect 259564 138892 259565 138956
rect 259499 138891 259565 138892
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 261342 97613 261402 139707
rect 262794 120454 263414 155898
rect 263550 142221 263610 188395
rect 263734 163437 263794 192475
rect 265022 168197 265082 204851
rect 266307 200836 266373 200837
rect 266307 200772 266308 200836
rect 266372 200772 266373 200836
rect 266307 200771 266373 200772
rect 265203 182884 265269 182885
rect 265203 182820 265204 182884
rect 265268 182820 265269 182884
rect 265203 182819 265269 182820
rect 265206 170917 265266 182819
rect 265203 170916 265269 170917
rect 265203 170852 265204 170916
rect 265268 170852 265269 170916
rect 265203 170851 265269 170852
rect 265019 168196 265085 168197
rect 265019 168132 265020 168196
rect 265084 168132 265085 168196
rect 265019 168131 265085 168132
rect 266310 164797 266370 200771
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 266307 164796 266373 164797
rect 266307 164732 266308 164796
rect 266372 164732 266373 164796
rect 266307 164731 266373 164732
rect 263731 163436 263797 163437
rect 263731 163372 263732 163436
rect 263796 163372 263797 163436
rect 263731 163371 263797 163372
rect 267294 160954 267914 196398
rect 271794 237454 272414 238000
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 269619 191180 269685 191181
rect 269619 191116 269620 191180
rect 269684 191116 269685 191180
rect 269619 191115 269685 191116
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 263547 142220 263613 142221
rect 263547 142156 263548 142220
rect 263612 142156 263613 142220
rect 263547 142155 263613 142156
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 261339 97612 261405 97613
rect 261339 97548 261340 97612
rect 261404 97548 261405 97612
rect 261339 97547 261405 97548
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 269622 3365 269682 191115
rect 271091 188596 271157 188597
rect 271091 188532 271092 188596
rect 271156 188532 271157 188596
rect 271091 188531 271157 188532
rect 271094 4045 271154 188531
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 276294 205954 276914 238000
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 275139 113524 275205 113525
rect 275139 113460 275140 113524
rect 275204 113460 275205 113524
rect 275139 113459 275205 113460
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271091 4044 271157 4045
rect 271091 3980 271092 4044
rect 271156 3980 271157 4044
rect 271091 3979 271157 3980
rect 269619 3364 269685 3365
rect 269619 3300 269620 3364
rect 269684 3300 269685 3364
rect 269619 3299 269685 3300
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 -4186 272414 20898
rect 275142 18597 275202 113459
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 275139 18596 275205 18597
rect 275139 18532 275140 18596
rect 275204 18532 275205 18596
rect 275139 18531 275205 18532
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 238000
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 238000
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 238000
rect 293174 235381 293234 309027
rect 293910 305421 293970 357307
rect 294294 357154 294914 367398
rect 293907 305420 293973 305421
rect 293907 305356 293908 305420
rect 293972 305356 293973 305420
rect 293907 305355 293973 305356
rect 295014 248301 295074 375259
rect 295382 312221 295442 578851
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 295563 367708 295629 367709
rect 295563 367644 295564 367708
rect 295628 367644 295629 367708
rect 295563 367643 295629 367644
rect 295379 312220 295445 312221
rect 295379 312156 295380 312220
rect 295444 312156 295445 312220
rect 295379 312155 295445 312156
rect 295379 257140 295445 257141
rect 295379 257076 295380 257140
rect 295444 257076 295445 257140
rect 295379 257075 295445 257076
rect 295011 248300 295077 248301
rect 295011 248236 295012 248300
rect 295076 248236 295077 248300
rect 295011 248235 295077 248236
rect 295382 240141 295442 257075
rect 295566 246261 295626 367643
rect 296483 358868 296549 358869
rect 296483 358804 296484 358868
rect 296548 358804 296549 358868
rect 296483 358803 296549 358804
rect 295563 246260 295629 246261
rect 295563 246196 295564 246260
rect 295628 246196 295629 246260
rect 295563 246195 295629 246196
rect 295379 240140 295445 240141
rect 295379 240076 295380 240140
rect 295444 240076 295445 240140
rect 295379 240075 295445 240076
rect 293171 235380 293237 235381
rect 293171 235316 293172 235380
rect 293236 235316 293237 235380
rect 293171 235315 293237 235316
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 294294 223954 294914 238000
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 291699 130116 291765 130117
rect 291699 130052 291700 130116
rect 291764 130052 291765 130116
rect 291699 130051 291765 130052
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 291702 58581 291762 130051
rect 293171 125900 293237 125901
rect 293171 125836 293172 125900
rect 293236 125836 293237 125900
rect 293171 125835 293237 125836
rect 293174 59941 293234 125835
rect 294294 115954 294914 151398
rect 295931 117604 295997 117605
rect 295931 117540 295932 117604
rect 295996 117540 295997 117604
rect 295931 117539 295997 117540
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 293171 59940 293237 59941
rect 293171 59876 293172 59940
rect 293236 59876 293237 59940
rect 293171 59875 293237 59876
rect 291699 58580 291765 58581
rect 291699 58516 291700 58580
rect 291764 58516 291765 58580
rect 291699 58515 291765 58516
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 295934 26893 295994 117539
rect 295931 26892 295997 26893
rect 295931 26828 295932 26892
rect 295996 26828 295997 26892
rect 295931 26827 295997 26828
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 296486 4045 296546 358803
rect 298507 357644 298573 357645
rect 298507 357580 298508 357644
rect 298572 357580 298573 357644
rect 298507 357579 298573 357580
rect 298510 240821 298570 357579
rect 298794 336454 299414 371898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 299979 359004 300045 359005
rect 299979 358940 299980 359004
rect 300044 358940 300045 359004
rect 299979 358939 300045 358940
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298507 240820 298573 240821
rect 298507 240756 298508 240820
rect 298572 240756 298573 240820
rect 298507 240755 298573 240756
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 296483 4044 296549 4045
rect 296483 3980 296484 4044
rect 296548 3980 296549 4044
rect 296483 3979 296549 3980
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 -2266 299414 11898
rect 299982 3501 300042 358939
rect 301451 356420 301517 356421
rect 301451 356356 301452 356420
rect 301516 356356 301517 356420
rect 301451 356355 301517 356356
rect 300163 135284 300229 135285
rect 300163 135220 300164 135284
rect 300228 135220 300229 135284
rect 300163 135219 300229 135220
rect 300166 69597 300226 135219
rect 300163 69596 300229 69597
rect 300163 69532 300164 69596
rect 300228 69532 300229 69596
rect 300163 69531 300229 69532
rect 301454 3637 301514 356355
rect 303294 340954 303914 376398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 304211 356284 304277 356285
rect 304211 356220 304212 356284
rect 304276 356220 304277 356284
rect 304211 356219 304277 356220
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 302739 101148 302805 101149
rect 302739 101084 302740 101148
rect 302804 101084 302805 101148
rect 302739 101083 302805 101084
rect 301635 100060 301701 100061
rect 301635 99996 301636 100060
rect 301700 99996 301701 100060
rect 301635 99995 301701 99996
rect 301638 62797 301698 99995
rect 301635 62796 301701 62797
rect 301635 62732 301636 62796
rect 301700 62732 301701 62796
rect 301635 62731 301701 62732
rect 302742 48925 302802 101083
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 302739 48924 302805 48925
rect 302739 48860 302740 48924
rect 302804 48860 302805 48924
rect 302739 48859 302805 48860
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 301451 3636 301517 3637
rect 301451 3572 301452 3636
rect 301516 3572 301517 3636
rect 301451 3571 301517 3572
rect 299979 3500 300045 3501
rect 299979 3436 299980 3500
rect 300044 3436 300045 3500
rect 299979 3435 300045 3436
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 -3226 303914 16398
rect 304214 4045 304274 356219
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 178000 308414 200898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 178000 312914 205398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 178000 317414 209898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 318011 186964 318077 186965
rect 318011 186900 318012 186964
rect 318076 186900 318077 186964
rect 318011 186899 318077 186900
rect 318014 177581 318074 186899
rect 320219 185604 320285 185605
rect 320219 185540 320220 185604
rect 320284 185540 320285 185604
rect 320219 185539 320285 185540
rect 318011 177580 318077 177581
rect 318011 177516 318012 177580
rect 318076 177516 318077 177580
rect 318011 177515 318077 177516
rect 306971 175676 307037 175677
rect 306971 175612 306972 175676
rect 307036 175612 307037 175676
rect 306971 175611 307037 175612
rect 306974 140045 307034 175611
rect 320222 171150 320282 185539
rect 321294 178954 321914 214398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 328499 467940 328565 467941
rect 328499 467876 328500 467940
rect 328564 467876 328565 467940
rect 328499 467875 328565 467876
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 327027 219332 327093 219333
rect 327027 219268 327028 219332
rect 327092 219268 327093 219332
rect 327027 219267 327093 219268
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 322059 181388 322125 181389
rect 322059 181324 322060 181388
rect 322124 181324 322125 181388
rect 322059 181323 322125 181324
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 178000 321914 178398
rect 321507 176220 321573 176221
rect 321507 176156 321508 176220
rect 321572 176156 321573 176220
rect 321507 176155 321573 176156
rect 321510 172141 321570 176155
rect 321507 172140 321573 172141
rect 321507 172076 321508 172140
rect 321572 172076 321573 172140
rect 321507 172075 321573 172076
rect 320222 171090 321386 171150
rect 321326 169829 321386 171090
rect 321323 169828 321389 169829
rect 321323 169764 321324 169828
rect 321388 169764 321389 169828
rect 321323 169763 321389 169764
rect 314208 151954 314528 151986
rect 314208 151718 314250 151954
rect 314486 151718 314528 151954
rect 314208 151634 314528 151718
rect 314208 151398 314250 151634
rect 314486 151398 314528 151634
rect 314208 151366 314528 151398
rect 317472 151954 317792 151986
rect 317472 151718 317514 151954
rect 317750 151718 317792 151954
rect 317472 151634 317792 151718
rect 317472 151398 317514 151634
rect 317750 151398 317792 151634
rect 317472 151366 317792 151398
rect 322062 150381 322122 181323
rect 322059 150380 322125 150381
rect 322059 150316 322060 150380
rect 322124 150316 322125 150380
rect 322059 150315 322125 150316
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 306971 140044 307037 140045
rect 306971 139980 306972 140044
rect 307036 139980 307037 140044
rect 306971 139979 307037 139980
rect 305499 139500 305565 139501
rect 305499 139436 305500 139500
rect 305564 139436 305565 139500
rect 305499 139435 305565 139436
rect 305502 37909 305562 139435
rect 307155 128076 307221 128077
rect 307155 128012 307156 128076
rect 307220 128012 307221 128076
rect 307155 128011 307221 128012
rect 305683 101284 305749 101285
rect 305683 101220 305684 101284
rect 305748 101220 305749 101284
rect 305683 101219 305749 101220
rect 305499 37908 305565 37909
rect 305499 37844 305500 37908
rect 305564 37844 305565 37908
rect 305499 37843 305565 37844
rect 305686 13021 305746 101219
rect 306971 97068 307037 97069
rect 306971 97004 306972 97068
rect 307036 97004 307037 97068
rect 306971 97003 307037 97004
rect 305683 13020 305749 13021
rect 305683 12956 305684 13020
rect 305748 12956 305749 13020
rect 305683 12955 305749 12956
rect 306974 8941 307034 97003
rect 307158 89181 307218 128011
rect 314208 115954 314528 115986
rect 314208 115718 314250 115954
rect 314486 115718 314528 115954
rect 314208 115634 314528 115718
rect 314208 115398 314250 115634
rect 314486 115398 314528 115634
rect 314208 115366 314528 115398
rect 317472 115954 317792 115986
rect 317472 115718 317514 115954
rect 317750 115718 317792 115954
rect 317472 115634 317792 115718
rect 317472 115398 317514 115634
rect 317750 115398 317792 115634
rect 317472 115366 317792 115398
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 325794 111454 326414 146898
rect 327030 139365 327090 219267
rect 327579 196756 327645 196757
rect 327579 196692 327580 196756
rect 327644 196692 327645 196756
rect 327579 196691 327645 196692
rect 327027 139364 327093 139365
rect 327027 139300 327028 139364
rect 327092 139300 327093 139364
rect 327027 139299 327093 139300
rect 327582 132157 327642 196691
rect 328502 142085 328562 467875
rect 330294 439954 330914 475398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 331259 452708 331325 452709
rect 331259 452644 331260 452708
rect 331324 452644 331325 452708
rect 331259 452643 331325 452644
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 328683 227764 328749 227765
rect 328683 227700 328684 227764
rect 328748 227700 328749 227764
rect 328683 227699 328749 227700
rect 328686 142221 328746 227699
rect 330294 223954 330914 259398
rect 331262 228989 331322 452643
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 332547 365804 332613 365805
rect 332547 365740 332548 365804
rect 332612 365740 332613 365804
rect 332547 365739 332613 365740
rect 331259 228988 331325 228989
rect 331259 228924 331260 228988
rect 331324 228924 331325 228988
rect 331259 228923 331325 228924
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 329787 220828 329853 220829
rect 329787 220764 329788 220828
rect 329852 220764 329853 220828
rect 329787 220763 329853 220764
rect 329790 143581 329850 220763
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 329787 143580 329853 143581
rect 329787 143516 329788 143580
rect 329852 143516 329853 143580
rect 329787 143515 329853 143516
rect 328683 142220 328749 142221
rect 328683 142156 328684 142220
rect 328748 142156 328749 142220
rect 328683 142155 328749 142156
rect 328499 142084 328565 142085
rect 328499 142020 328500 142084
rect 328564 142020 328565 142084
rect 328499 142019 328565 142020
rect 327579 132156 327645 132157
rect 327579 132092 327580 132156
rect 327644 132092 327645 132156
rect 327579 132091 327645 132092
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307155 89180 307221 89181
rect 307155 89116 307156 89180
rect 307220 89116 307221 89180
rect 307155 89115 307221 89116
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 306971 8940 307037 8941
rect 306971 8876 306972 8940
rect 307036 8876 307037 8940
rect 306971 8875 307037 8876
rect 304211 4044 304277 4045
rect 304211 3980 304212 4044
rect 304276 3980 304277 4044
rect 304211 3979 304277 3980
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 61954 312914 94000
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 66454 317414 94000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 70954 321914 94000
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 115954 330914 151398
rect 331262 131749 331322 228923
rect 331259 131748 331325 131749
rect 331259 131684 331260 131748
rect 331324 131684 331325 131748
rect 331259 131683 331325 131684
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 332550 3501 332610 365739
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 340827 360228 340893 360229
rect 340827 360164 340828 360228
rect 340892 360164 340893 360228
rect 340827 360163 340893 360164
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 338251 223684 338317 223685
rect 338251 223620 338252 223684
rect 338316 223620 338317 223684
rect 338251 223619 338317 223620
rect 336779 213212 336845 213213
rect 336779 213148 336780 213212
rect 336844 213148 336845 213212
rect 336779 213147 336845 213148
rect 335675 195260 335741 195261
rect 335675 195196 335676 195260
rect 335740 195196 335741 195260
rect 335675 195195 335741 195196
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 332731 178668 332797 178669
rect 332731 178604 332732 178668
rect 332796 178604 332797 178668
rect 332731 178603 332797 178604
rect 332734 123317 332794 178603
rect 334019 177444 334085 177445
rect 334019 177380 334020 177444
rect 334084 177380 334085 177444
rect 334019 177379 334085 177380
rect 334022 165749 334082 177379
rect 334019 165748 334085 165749
rect 334019 165684 334020 165748
rect 334084 165684 334085 165748
rect 334019 165683 334085 165684
rect 334794 156454 335414 191898
rect 335678 180810 335738 195195
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 332731 123316 332797 123317
rect 332731 123252 332732 123316
rect 332796 123252 332797 123316
rect 332731 123251 332797 123252
rect 334794 120454 335414 155898
rect 335494 180750 335738 180810
rect 335494 132510 335554 180750
rect 335675 180164 335741 180165
rect 335675 180100 335676 180164
rect 335740 180100 335741 180164
rect 335675 180099 335741 180100
rect 335678 160173 335738 180099
rect 335675 160172 335741 160173
rect 335675 160108 335676 160172
rect 335740 160108 335741 160172
rect 335675 160107 335741 160108
rect 335494 132450 335738 132510
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 335678 116109 335738 132450
rect 335675 116108 335741 116109
rect 335675 116044 335676 116108
rect 335740 116044 335741 116108
rect 335675 116043 335741 116044
rect 336782 109173 336842 213147
rect 336963 177308 337029 177309
rect 336963 177244 336964 177308
rect 337028 177244 337029 177308
rect 336963 177243 337029 177244
rect 336966 140861 337026 177243
rect 336963 140860 337029 140861
rect 336963 140796 336964 140860
rect 337028 140796 337029 140860
rect 336963 140795 337029 140796
rect 338254 115973 338314 223619
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 338251 115972 338317 115973
rect 338251 115908 338252 115972
rect 338316 115908 338317 115972
rect 338251 115907 338317 115908
rect 336779 109172 336845 109173
rect 336779 109108 336780 109172
rect 336844 109108 336845 109172
rect 336779 109107 336845 109108
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 332547 3500 332613 3501
rect 332547 3436 332548 3500
rect 332612 3436 332613 3500
rect 332547 3435 332613 3436
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 340830 3501 340890 360163
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 342299 179212 342365 179213
rect 342299 179148 342300 179212
rect 342364 179148 342365 179212
rect 342299 179147 342365 179148
rect 342302 135285 342362 179147
rect 343794 165454 344414 200898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 345059 196620 345125 196621
rect 345059 196556 345060 196620
rect 345124 196556 345125 196620
rect 345059 196555 345125 196556
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 342299 135284 342365 135285
rect 342299 135220 342300 135284
rect 342364 135220 342365 135284
rect 342299 135219 342365 135220
rect 343794 129454 344414 164898
rect 345062 161533 345122 196555
rect 346347 179348 346413 179349
rect 346347 179284 346348 179348
rect 346412 179284 346413 179348
rect 346347 179283 346413 179284
rect 345059 161532 345125 161533
rect 345059 161468 345060 161532
rect 345124 161468 345125 161532
rect 345059 161467 345125 161468
rect 346350 139501 346410 179283
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 346347 139500 346413 139501
rect 346347 139436 346348 139500
rect 346412 139436 346413 139500
rect 346347 139435 346413 139436
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 340827 3500 340893 3501
rect 340827 3436 340828 3500
rect 340892 3436 340893 3500
rect 340827 3435 340893 3436
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< obsm4 >>
rect 68800 174494 96960 174600
rect 97020 174494 98320 174600
rect 98380 174494 99408 174600
rect 99468 174494 100768 174600
rect 100828 174494 101992 174600
rect 102052 174494 103352 174600
rect 103412 174494 104576 174600
rect 104636 174494 105664 174600
rect 105724 174494 107024 174600
rect 107084 174494 108112 174600
rect 108172 174494 109472 174600
rect 109532 174494 110696 174600
rect 110756 174494 112056 174600
rect 112116 174494 113144 174600
rect 113204 174494 114368 174600
rect 114428 174494 115728 174600
rect 115788 174494 116952 174600
rect 117012 174494 118312 174600
rect 118372 174494 119400 174600
rect 119460 174494 120760 174600
rect 120820 174494 121848 174600
rect 121908 174494 123072 174600
rect 123132 174494 124432 174600
rect 124492 174494 125656 174600
rect 125716 174494 127016 174600
rect 127076 174494 128104 174600
rect 128164 174494 129464 174600
rect 129524 174494 130688 174600
rect 130748 174494 132048 174600
rect 132108 174494 133136 174600
rect 133196 174494 134360 174600
rect 134420 174494 135720 174600
rect 135780 174494 148232 174600
rect 148292 174494 158840 174600
rect 158900 174494 164756 174600
rect 68800 151986 164756 174494
rect 68800 151366 69072 151986
rect 69420 151366 164136 151986
rect 164484 151366 164756 151986
rect 68800 147486 164756 151366
rect 68800 146866 69752 147486
rect 70100 146866 163456 147486
rect 163804 146866 164756 147486
rect 68800 115986 164756 146866
rect 68800 115366 69072 115986
rect 69420 115366 164136 115986
rect 164484 115366 164756 115986
rect 68800 111486 164756 115366
rect 68800 110866 69752 111486
rect 70100 110866 163456 111486
rect 163804 110866 164756 111486
rect 68800 95200 164756 110866
rect 68800 95100 74656 95200
rect 74716 95100 84312 95200
rect 84372 95100 85536 95200
rect 85596 95100 86624 95200
rect 86684 95100 87984 95200
rect 88044 95100 88936 95200
rect 88996 95100 90160 95200
rect 90220 95100 91384 95200
rect 91444 95100 92472 95200
rect 92532 95100 93832 95200
rect 93892 95100 94920 95200
rect 94980 95100 96008 95200
rect 96068 95100 96688 95200
rect 96748 95100 97096 95200
rect 97156 95100 98048 95200
rect 98108 95100 98456 95200
rect 98516 95100 99136 95200
rect 99196 95100 99544 95200
rect 99604 95100 100632 95200
rect 100692 95100 100768 95200
rect 100828 95100 101856 95200
rect 101916 95100 101992 95200
rect 102052 95100 102944 95200
rect 103004 95100 103216 95200
rect 103276 95100 104304 95200
rect 104364 95100 104440 95200
rect 104500 95100 105392 95200
rect 105452 95100 105664 95200
rect 105724 95100 106480 95200
rect 106540 95100 106616 95200
rect 106676 95100 107704 95200
rect 107764 95100 108112 95200
rect 108172 95100 109064 95200
rect 109124 95100 109472 95200
rect 109532 95100 110152 95200
rect 110212 95100 110696 95200
rect 110756 95100 111240 95200
rect 111300 95100 111920 95200
rect 111980 95100 112328 95200
rect 112388 95100 113144 95200
rect 113204 95100 113688 95200
rect 113748 95100 114368 95200
rect 114428 95100 114776 95200
rect 114836 95100 115456 95200
rect 115516 95100 115864 95200
rect 115924 95100 116680 95200
rect 116740 95100 117088 95200
rect 117148 95100 117904 95200
rect 117964 95100 118176 95200
rect 118236 95100 119400 95200
rect 119460 95100 119536 95200
rect 119596 95100 120216 95200
rect 120276 95100 120624 95200
rect 120684 95100 121712 95200
rect 121772 95100 121984 95200
rect 122044 95100 122800 95200
rect 122860 95100 123208 95200
rect 123268 95100 124024 95200
rect 124084 95100 124432 95200
rect 124492 95100 125384 95200
rect 125444 95100 125656 95200
rect 125716 95100 126472 95200
rect 126532 95100 126608 95200
rect 126668 95100 128104 95200
rect 128164 95100 129328 95200
rect 129388 95100 130688 95200
rect 130748 95100 131912 95200
rect 131972 95100 133136 95200
rect 133196 95100 134360 95200
rect 134420 95100 135584 95200
rect 135644 95100 151496 95200
rect 151556 95100 151632 95200
rect 151692 95100 151768 95200
rect 151828 95100 151904 95200
rect 151964 95100 164756 95200
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 68250 579218 68486 579454
rect 68250 578898 68486 579134
rect 98970 579218 99206 579454
rect 98970 578898 99206 579134
rect 129690 579218 129926 579454
rect 129690 578898 129926 579134
rect 160410 579218 160646 579454
rect 160410 578898 160646 579134
rect 191130 579218 191366 579454
rect 191130 578898 191366 579134
rect 221850 579218 222086 579454
rect 221850 578898 222086 579134
rect 83610 547718 83846 547954
rect 83610 547398 83846 547634
rect 114330 547718 114566 547954
rect 114330 547398 114566 547634
rect 145050 547718 145286 547954
rect 145050 547398 145286 547634
rect 175770 547718 176006 547954
rect 175770 547398 176006 547634
rect 206490 547718 206726 547954
rect 206490 547398 206726 547634
rect 237210 547718 237446 547954
rect 237210 547398 237446 547634
rect 68250 543218 68486 543454
rect 68250 542898 68486 543134
rect 98970 543218 99206 543454
rect 98970 542898 99206 543134
rect 129690 543218 129926 543454
rect 129690 542898 129926 543134
rect 160410 543218 160646 543454
rect 160410 542898 160646 543134
rect 191130 543218 191366 543454
rect 191130 542898 191366 543134
rect 221850 543218 222086 543454
rect 221850 542898 222086 543134
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 83610 511718 83846 511954
rect 83610 511398 83846 511634
rect 114330 511718 114566 511954
rect 114330 511398 114566 511634
rect 145050 511718 145286 511954
rect 145050 511398 145286 511634
rect 175770 511718 176006 511954
rect 175770 511398 176006 511634
rect 206490 511718 206726 511954
rect 206490 511398 206726 511634
rect 237210 511718 237446 511954
rect 237210 511398 237446 511634
rect 68250 507218 68486 507454
rect 68250 506898 68486 507134
rect 98970 507218 99206 507454
rect 98970 506898 99206 507134
rect 129690 507218 129926 507454
rect 129690 506898 129926 507134
rect 160410 507218 160646 507454
rect 160410 506898 160646 507134
rect 191130 507218 191366 507454
rect 191130 506898 191366 507134
rect 221850 507218 222086 507454
rect 221850 506898 222086 507134
rect 83610 475718 83846 475954
rect 83610 475398 83846 475634
rect 114330 475718 114566 475954
rect 114330 475398 114566 475634
rect 145050 475718 145286 475954
rect 145050 475398 145286 475634
rect 175770 475718 176006 475954
rect 175770 475398 176006 475634
rect 206490 475718 206726 475954
rect 206490 475398 206726 475634
rect 237210 475718 237446 475954
rect 237210 475398 237446 475634
rect 68250 471218 68486 471454
rect 68250 470898 68486 471134
rect 98970 471218 99206 471454
rect 98970 470898 99206 471134
rect 129690 471218 129926 471454
rect 129690 470898 129926 471134
rect 160410 471218 160646 471454
rect 160410 470898 160646 471134
rect 191130 471218 191366 471454
rect 191130 470898 191366 471134
rect 221850 471218 222086 471454
rect 221850 470898 222086 471134
rect 83610 439718 83846 439954
rect 83610 439398 83846 439634
rect 114330 439718 114566 439954
rect 114330 439398 114566 439634
rect 145050 439718 145286 439954
rect 145050 439398 145286 439634
rect 175770 439718 176006 439954
rect 175770 439398 176006 439634
rect 206490 439718 206726 439954
rect 206490 439398 206726 439634
rect 237210 439718 237446 439954
rect 237210 439398 237446 439634
rect 68250 435218 68486 435454
rect 68250 434898 68486 435134
rect 98970 435218 99206 435454
rect 98970 434898 99206 435134
rect 129690 435218 129926 435454
rect 129690 434898 129926 435134
rect 160410 435218 160646 435454
rect 160410 434898 160646 435134
rect 191130 435218 191366 435454
rect 191130 434898 191366 435134
rect 221850 435218 222086 435454
rect 221850 434898 222086 435134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 89610 259718 89846 259954
rect 89610 259398 89846 259634
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 69128 151718 69364 151954
rect 69128 151398 69364 151634
rect 164192 151718 164428 151954
rect 164192 151398 164428 151634
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 115718 69364 115954
rect 69128 115398 69364 115634
rect 164192 115718 164428 115954
rect 164192 115398 164428 115634
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 199610 331718 199846 331954
rect 199610 331398 199846 331634
rect 230330 331718 230566 331954
rect 230330 331398 230566 331634
rect 261050 331718 261286 331954
rect 261050 331398 261286 331634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 184250 327218 184486 327454
rect 184250 326898 184486 327134
rect 214970 327218 215206 327454
rect 214970 326898 215206 327134
rect 245690 327218 245926 327454
rect 245690 326898 245926 327134
rect 276410 327218 276646 327454
rect 276410 326898 276646 327134
rect 199610 295718 199846 295954
rect 199610 295398 199846 295634
rect 230330 295718 230566 295954
rect 230330 295398 230566 295634
rect 261050 295718 261286 295954
rect 261050 295398 261286 295634
rect 184250 291218 184486 291454
rect 184250 290898 184486 291134
rect 214970 291218 215206 291454
rect 214970 290898 215206 291134
rect 245690 291218 245926 291454
rect 245690 290898 245926 291134
rect 276410 291218 276646 291454
rect 276410 290898 276646 291134
rect 199610 259718 199846 259954
rect 199610 259398 199846 259634
rect 230330 259718 230566 259954
rect 230330 259398 230566 259634
rect 261050 259718 261286 259954
rect 261050 259398 261286 259634
rect 184250 255218 184486 255454
rect 184250 254898 184486 255134
rect 214970 255218 215206 255454
rect 214970 254898 215206 255134
rect 245690 255218 245926 255454
rect 245690 254898 245926 255134
rect 276410 255218 276646 255454
rect 276410 254898 276646 255134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 227916 151718 228152 151954
rect 227916 151398 228152 151634
rect 237847 151718 238083 151954
rect 237847 151398 238083 151634
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 227916 115718 228152 115954
rect 227916 115398 228152 115634
rect 237847 115718 238083 115954
rect 237847 115398 238083 115634
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 242813 110898 243049 111134
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 314250 151718 314486 151954
rect 314250 151398 314486 151634
rect 317514 151718 317750 151954
rect 317514 151398 317750 151634
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 314250 115718 314486 115954
rect 314250 115398 314486 115634
rect 317514 115718 317750 115954
rect 317514 115398 317750 115634
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 68250 579454
rect 68486 579218 98970 579454
rect 99206 579218 129690 579454
rect 129926 579218 160410 579454
rect 160646 579218 191130 579454
rect 191366 579218 221850 579454
rect 222086 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 68250 579134
rect 68486 578898 98970 579134
rect 99206 578898 129690 579134
rect 129926 578898 160410 579134
rect 160646 578898 191130 579134
rect 191366 578898 221850 579134
rect 222086 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 83610 547954
rect 83846 547718 114330 547954
rect 114566 547718 145050 547954
rect 145286 547718 175770 547954
rect 176006 547718 206490 547954
rect 206726 547718 237210 547954
rect 237446 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 83610 547634
rect 83846 547398 114330 547634
rect 114566 547398 145050 547634
rect 145286 547398 175770 547634
rect 176006 547398 206490 547634
rect 206726 547398 237210 547634
rect 237446 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 68250 543454
rect 68486 543218 98970 543454
rect 99206 543218 129690 543454
rect 129926 543218 160410 543454
rect 160646 543218 191130 543454
rect 191366 543218 221850 543454
rect 222086 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 68250 543134
rect 68486 542898 98970 543134
rect 99206 542898 129690 543134
rect 129926 542898 160410 543134
rect 160646 542898 191130 543134
rect 191366 542898 221850 543134
rect 222086 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 83610 511954
rect 83846 511718 114330 511954
rect 114566 511718 145050 511954
rect 145286 511718 175770 511954
rect 176006 511718 206490 511954
rect 206726 511718 237210 511954
rect 237446 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 83610 511634
rect 83846 511398 114330 511634
rect 114566 511398 145050 511634
rect 145286 511398 175770 511634
rect 176006 511398 206490 511634
rect 206726 511398 237210 511634
rect 237446 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 68250 507454
rect 68486 507218 98970 507454
rect 99206 507218 129690 507454
rect 129926 507218 160410 507454
rect 160646 507218 191130 507454
rect 191366 507218 221850 507454
rect 222086 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 68250 507134
rect 68486 506898 98970 507134
rect 99206 506898 129690 507134
rect 129926 506898 160410 507134
rect 160646 506898 191130 507134
rect 191366 506898 221850 507134
rect 222086 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 83610 475954
rect 83846 475718 114330 475954
rect 114566 475718 145050 475954
rect 145286 475718 175770 475954
rect 176006 475718 206490 475954
rect 206726 475718 237210 475954
rect 237446 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 83610 475634
rect 83846 475398 114330 475634
rect 114566 475398 145050 475634
rect 145286 475398 175770 475634
rect 176006 475398 206490 475634
rect 206726 475398 237210 475634
rect 237446 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 68250 471454
rect 68486 471218 98970 471454
rect 99206 471218 129690 471454
rect 129926 471218 160410 471454
rect 160646 471218 191130 471454
rect 191366 471218 221850 471454
rect 222086 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 68250 471134
rect 68486 470898 98970 471134
rect 99206 470898 129690 471134
rect 129926 470898 160410 471134
rect 160646 470898 191130 471134
rect 191366 470898 221850 471134
rect 222086 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 83610 439954
rect 83846 439718 114330 439954
rect 114566 439718 145050 439954
rect 145286 439718 175770 439954
rect 176006 439718 206490 439954
rect 206726 439718 237210 439954
rect 237446 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 83610 439634
rect 83846 439398 114330 439634
rect 114566 439398 145050 439634
rect 145286 439398 175770 439634
rect 176006 439398 206490 439634
rect 206726 439398 237210 439634
rect 237446 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 68250 435454
rect 68486 435218 98970 435454
rect 99206 435218 129690 435454
rect 129926 435218 160410 435454
rect 160646 435218 191130 435454
rect 191366 435218 221850 435454
rect 222086 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 68250 435134
rect 68486 434898 98970 435134
rect 99206 434898 129690 435134
rect 129926 434898 160410 435134
rect 160646 434898 191130 435134
rect 191366 434898 221850 435134
rect 222086 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 199610 331954
rect 199846 331718 230330 331954
rect 230566 331718 261050 331954
rect 261286 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 199610 331634
rect 199846 331398 230330 331634
rect 230566 331398 261050 331634
rect 261286 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 184250 327454
rect 184486 327218 214970 327454
rect 215206 327218 245690 327454
rect 245926 327218 276410 327454
rect 276646 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 184250 327134
rect 184486 326898 214970 327134
rect 215206 326898 245690 327134
rect 245926 326898 276410 327134
rect 276646 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 199610 295954
rect 199846 295718 230330 295954
rect 230566 295718 261050 295954
rect 261286 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 199610 295634
rect 199846 295398 230330 295634
rect 230566 295398 261050 295634
rect 261286 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 184250 291454
rect 184486 291218 214970 291454
rect 215206 291218 245690 291454
rect 245926 291218 276410 291454
rect 276646 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 184250 291134
rect 184486 290898 214970 291134
rect 215206 290898 245690 291134
rect 245926 290898 276410 291134
rect 276646 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 89610 259954
rect 89846 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 199610 259954
rect 199846 259718 230330 259954
rect 230566 259718 261050 259954
rect 261286 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 89610 259634
rect 89846 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 199610 259634
rect 199846 259398 230330 259634
rect 230566 259398 261050 259634
rect 261286 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 184250 255454
rect 184486 255218 214970 255454
rect 215206 255218 245690 255454
rect 245926 255218 276410 255454
rect 276646 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 184250 255134
rect 184486 254898 214970 255134
rect 215206 254898 245690 255134
rect 245926 254898 276410 255134
rect 276646 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 69128 151954
rect 69364 151718 164192 151954
rect 164428 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 227916 151954
rect 228152 151718 237847 151954
rect 238083 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 314250 151954
rect 314486 151718 317514 151954
rect 317750 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 69128 151634
rect 69364 151398 164192 151634
rect 164428 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 227916 151634
rect 228152 151398 237847 151634
rect 238083 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 314250 151634
rect 314486 151398 317514 151634
rect 317750 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 69128 115954
rect 69364 115718 164192 115954
rect 164428 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 227916 115954
rect 228152 115718 237847 115954
rect 238083 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 314250 115954
rect 314486 115718 317514 115954
rect 317750 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 69128 115634
rect 69364 115398 164192 115634
rect 164428 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 227916 115634
rect 228152 115398 237847 115634
rect 238083 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 314250 115634
rect 314486 115398 317514 115634
rect 317750 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_etpu  wrapped_etpu_3
timestamp 0
transform 1 0 64000 0 1 405000
box -10 0 180000 180000
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
use wrapped_ibnalhaytham  wrapped_ibnalhaytham_1
timestamp 0
transform 1 0 180000 0 1 240000
box 0 0 113010 115154
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 176600 74414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 294000 74414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 587000 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 176600 110414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 294000 110414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 587000 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 176600 146414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 587000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 357154 182414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 587000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 178000 218414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 357154 218414 403000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 587000 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 357154 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 357154 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 176600 83414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 294000 83414 403000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 587000 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 176600 119414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 294000 119414 403000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 587000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 176600 155414 403000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 587000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 587000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 178000 227414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 587000 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 357154 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 176600 92414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 294000 92414 403000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 587000 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 176600 128414 403000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 587000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 176600 164414 403000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 587000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 587000 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 178000 236414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 587000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 357154 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 178000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 403000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 587000 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 294000 101414 403000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 587000 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 176600 137414 403000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 587000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 403000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 587000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 587000 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 587000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 357154 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 178000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 294000 96914 403000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 587000 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 176600 132914 403000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 587000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 403000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 587000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 587000 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 587000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 357154 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 178000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 176600 69914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 294000 69914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 587000 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 176600 105914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 294000 105914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 587000 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 176600 141914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 587000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 587000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 357154 213914 403000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 587000 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 178000 249914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 357154 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 357154 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 178000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 176600 78914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 294000 78914 403000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 587000 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 176600 114914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 294000 114914 403000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 587000 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 176600 150914 403000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 587000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 587000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 178000 222914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 587000 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 357154 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 357154 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 176600 87914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 294000 87914 403000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 587000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 176600 123914 403000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 587000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 176600 159914 403000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 587000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 587000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 178000 231914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 587000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 357154 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
